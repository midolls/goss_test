magic
tech sky130A
magscale 1 2
timestamp 1691578050
<< metal1 >>
rect 1470 2726 1576 2790
rect 4304 2762 4504 2766
rect 4304 2678 4524 2762
rect 1590 2256 1696 2320
rect 2184 2252 2282 2280
rect 2184 2242 2298 2252
rect 2200 2214 2298 2242
rect 4322 2248 4358 2250
rect 4322 2214 4394 2248
rect 2052 2170 2116 2176
rect 2052 2118 2058 2170
rect 2110 2118 2116 2170
rect 2052 2112 2116 2118
rect 1480 1768 1588 1834
rect 2048 1376 2112 1382
rect 2048 1324 2054 1376
rect 2108 1366 2112 1376
rect 4354 1368 4394 2214
rect 2108 1330 2280 1366
rect 4322 1334 4394 1368
rect 4322 1332 4358 1334
rect 2108 1324 2112 1330
rect 2048 1318 2112 1324
rect 4426 904 4524 2678
rect 4304 816 4524 904
<< via1 >>
rect 2058 2118 2110 2170
rect 2054 1324 2108 1376
<< metal2 >>
rect 2052 2170 2116 2176
rect 2052 2118 2058 2170
rect 2110 2118 2116 2170
rect 2052 2112 2116 2118
rect 2058 1382 2106 2112
rect 2048 1376 2112 1382
rect 2048 1324 2054 1376
rect 2108 1324 2112 1376
rect 2048 1318 2112 1324
use nand  x1
timestamp 1691241966
transform 1 0 988 0 1 1958
box 478 -206 1312 848
use inverter  x2
timestamp 1691573807
transform 1 0 1966 0 1 1800
box 314 -10 738 970
use inverter  x3
timestamp 1691573807
transform 1 0 2373 0 1 1800
box 314 -10 738 970
use inverter  x4
timestamp 1691573807
transform 1 0 2778 0 1 1800
box 314 -10 738 970
use inverter  x5
timestamp 1691573807
transform 1 0 3182 0 1 1800
box 314 -10 738 970
use inverter  x6
timestamp 1691573807
transform 1 0 3588 0 1 1800
box 314 -10 738 970
use inverter  x7
timestamp 1691573807
transform -1 0 4640 0 -1 1782
box 314 -10 738 970
use inverter  x8
timestamp 1691573807
transform -1 0 4234 0 -1 1782
box 314 -10 738 970
use inverter  x9
timestamp 1691573807
transform -1 0 3830 0 -1 1782
box 314 -10 738 970
use inverter  x10
timestamp 1691573807
transform -1 0 3426 0 -1 1782
box 314 -10 738 970
use inverter  x11
timestamp 1691573807
transform -1 0 3018 0 -1 1782
box 314 -10 738 970
<< labels >>
flabel metal1 1470 2726 1576 2790 0 FreeSans 160 0 0 0 VDD
port 0 nsew
flabel metal1 1482 1770 1588 1834 0 FreeSans 160 0 0 0 VSS
port 1 nsew
flabel metal1 1590 2256 1696 2320 0 FreeSans 160 0 0 0 EN
port 3 nsew
flabel metal1 2154 1330 2250 1360 0 FreeSans 160 0 0 0 CLK
port 5 nsew
<< end >>
