magic
tech sky130A
magscale 1 2
timestamp 1690721753
<< error_p >>
rect -29 -95 29 -89
rect -29 -129 -17 -95
rect -29 -135 29 -129
<< nwell >>
rect -211 -268 211 268
<< pmos >>
rect -15 -48 15 120
<< pdiff >>
rect -73 108 -15 120
rect -73 -36 -61 108
rect -27 -36 -15 108
rect -73 -48 -15 -36
rect 15 108 73 120
rect 15 -36 27 108
rect 61 -36 73 108
rect 15 -48 73 -36
<< pdiffc >>
rect -61 -36 -27 108
rect 27 -36 61 108
<< nsubdiff >>
rect -175 198 -79 232
rect 79 198 175 232
rect -175 135 -141 198
rect 141 135 175 198
rect -175 -198 -141 -135
rect 141 -198 175 -135
rect -175 -232 -79 -198
rect 79 -232 175 -198
<< nsubdiffcont >>
rect -79 198 79 232
rect -175 -135 -141 135
rect 141 -135 175 135
rect -79 -232 79 -198
<< poly >>
rect -15 120 15 146
rect -15 -79 15 -48
rect -33 -95 33 -79
rect -33 -129 -17 -95
rect 17 -129 33 -95
rect -33 -145 33 -129
<< polycont >>
rect -17 -129 17 -95
<< locali >>
rect -175 198 -79 232
rect 79 198 175 232
rect -175 135 -141 198
rect 141 135 175 198
rect -61 108 -27 124
rect -61 -52 -27 -36
rect 27 108 61 124
rect 27 -52 61 -36
rect -33 -129 -17 -95
rect 17 -129 33 -95
rect -175 -198 -141 -135
rect 141 -198 175 -135
rect -175 -232 -79 -198
rect 79 -232 175 -198
<< viali >>
rect -61 -36 -27 108
rect 27 -36 61 108
rect -17 -129 17 -95
<< metal1 >>
rect -67 108 -21 120
rect -67 -36 -61 108
rect -27 -36 -21 108
rect -67 -48 -21 -36
rect 21 108 67 120
rect 21 -36 27 108
rect 61 -36 67 108
rect 21 -48 67 -36
rect -29 -95 29 -89
rect -29 -129 -17 -95
rect 17 -129 29 -95
rect -29 -135 29 -129
<< properties >>
string FIXED_BBOX -158 -215 158 215
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.84 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
