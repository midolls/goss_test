* NGSPICE file created from inverter.ext - technology: sky130A

.subckt inverter Vin Vout VDD VSS
X0 Vout.t0 Vin.t0 VSS.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1 Vout.t1 Vin.t1 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
R0 Vin.n0 Vin.t1 222.611
R1 Vin Vin.t0 140.625
R2 Vin.n0 Vin 0.6255
R3 Vin Vin.n0 0.038
R4 VSS.n9 VSS.n4 451.942
R5 VSS.n1 VSS.n0 390.688
R6 VSS.n3 VSS.n2 86.9652
R7 VSS.n15 VSS.n14 86.2123
R8 VSS.n12 VSS.t1 41.7354
R9 VSS.n10 VSS.n3 28.5262
R10 VSS.n16 VSS.n15 9.3005
R11 VSS.n9 VSS.n6 5.79462
R12 VSS.n6 VSS.n5 4.95547
R13 VSS.n11 VSS.n10 0.366214
R14 VSS.n10 VSS.n9 0.218539
R15 VSS.n9 VSS.t0 0.218539
R16 VSS VSS.n16 0.168867
R17 VSS.n8 VSS.n7 0.10956
R18 VSS.t0 VSS.n8 0.10956
R19 VSS.n14 VSS.n13 0.0944005
R20 VSS.n2 VSS.n1 0.0944005
R21 VSS.n12 VSS.n11 0.0630582
R22 VSS.n16 VSS.n12 0.0425918
R23 Vout Vout.t0 42.4673
R24 Vout Vout.t1 35.2375
R25 VDD.n3 VDD.n2 185
R26 VDD.n12 VDD.n11 185
R27 VDD.t0 VDD.n4 158.304
R28 VDD.t0 VDD.n7 158.304
R29 VDD.n12 VDD.n10 104.659
R30 VDD.n3 VDD.n1 104.659
R31 VDD.n14 VDD.t1 34.3985
R32 VDD.n13 VDD.n3 29.3652
R33 VDD.n13 VDD.n12 29.3652
R34 VDD VDD.n14 0.20675
R35 VDD.n14 VDD.n13 0.0598937
R36 VDD.n6 VDD.n5 0.0349892
R37 VDD.t0 VDD.n6 0.0349892
R38 VDD.n10 VDD.n9 0.018623
R39 VDD.n1 VDD.n0 0.018623
R40 VDD.n13 VDD.n8 0.00390556
R41 VDD.n8 VDD.t0 0.00390556
C0 Vout Vin 0.166f
C1 Vout VDD 0.326f
C2 Vin VDD 0.25f
.ends

