* NGSPICE file created from ringosil.ext - technology: sky130A

.subckt ringosil CLK EN_CLK VSS VDD
X0 x7.Vin x6.Vin VDD.t11 VDD.t10 sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X1 VDD.t13 x11.Vin CLK.t1 VDD.t12 sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X2 VSS.t16 x8.Vin x9.Vin VSS.t15 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X3 x4.Vin x3.Vin VSS.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X4 x5.Vin x4.Vin VSS.t7 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X5 x5.Vin x4.Vin VDD.t7 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X6 x6.Vin x5.Vin VDD.t21 VDD.t20 sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X7 VSS.t11 x11.Vin CLK.t0 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X8 VDD.t5 x9.Vout x11.Vin VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X9 x7.Vin x6.Vin VSS.t9 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X10 x3.Vin x2.Vin VDD.t23 VDD.t22 sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X11 x2.Vin EN_CLK.t0 VDD.t17 VDD.t16 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X12 a_1692_1940# EN_CLK.t1 VSS.t14 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X13 x6.Vin x5.Vin VSS.t17 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X14 VSS.t6 x9.Vout x11.Vin VSS.t5 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X15 VDD.t3 x9.Vin x9.Vout VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X16 x3.Vin x2.Vin VSS.t18 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X17 VDD.t15 x7.Vin x8.Vin VDD.t14 sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X18 VDD.t9 CLK.t2 x2.Vin VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X19 x2.Vin CLK.t3 a_1692_1940# VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X20 VSS.t3 x9.Vin x9.Vout VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X21 x4.Vin x3.Vin VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X22 VSS.t12 x7.Vin x8.Vin VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X23 VDD.t19 x8.Vin x9.Vin VDD.t18 sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
R0 VDD.n130 VDD.n129 4346.59
R1 VDD.n124 VDD.n8 1256.47
R2 VDD.n128 VDD.n8 1256.47
R3 VDD.n124 VDD.n9 1256.47
R4 VDD.n128 VDD.n9 1256.47
R5 VDD.n117 VDD.n11 1256.47
R6 VDD.n121 VDD.n11 1256.47
R7 VDD.n117 VDD.n12 1256.47
R8 VDD.n121 VDD.n12 1256.47
R9 VDD.n110 VDD.n14 1256.47
R10 VDD.n114 VDD.n14 1256.47
R11 VDD.n110 VDD.n15 1256.47
R12 VDD.n114 VDD.n15 1256.47
R13 VDD.n103 VDD.n17 1256.47
R14 VDD.n107 VDD.n17 1256.47
R15 VDD.n103 VDD.n18 1256.47
R16 VDD.n107 VDD.n18 1256.47
R17 VDD.n100 VDD.n20 1256.47
R18 VDD.n96 VDD.n21 1256.47
R19 VDD.n100 VDD.n21 1256.47
R20 VDD.n26 VDD.n25 1256.47
R21 VDD.n77 VDD.n25 1256.47
R22 VDD.n77 VDD.n23 1256.47
R23 VDD.n74 VDD.n28 1256.47
R24 VDD.n37 VDD.n28 1256.47
R25 VDD.n74 VDD.n29 1256.47
R26 VDD.n37 VDD.n29 1256.47
R27 VDD.n39 VDD.n36 1256.47
R28 VDD.n66 VDD.n36 1256.47
R29 VDD.n39 VDD.n34 1256.47
R30 VDD.n66 VDD.n34 1256.47
R31 VDD.n63 VDD.n41 1256.47
R32 VDD.n50 VDD.n41 1256.47
R33 VDD.n63 VDD.n42 1256.47
R34 VDD.n50 VDD.n42 1256.47
R35 VDD.n54 VDD.n48 1256.47
R36 VDD.n54 VDD.n49 1256.47
R37 VDD.n56 VDD.n48 1256.47
R38 VDD.n131 VDD.n5 1108.24
R39 VDD.n135 VDD.n5 1108.24
R40 VDD.n131 VDD.n6 1108.24
R41 VDD.n135 VDD.n6 1108.24
R42 VDD.n141 VDD.n3 1108.24
R43 VDD.n141 VDD.n4 1108.24
R44 VDD.n139 VDD.n3 1108.24
R45 VDD.n130 VDD.t8 332.08
R46 VDD.n136 VDD.t8 332.08
R47 VDD.t16 VDD.n137 332.08
R48 VDD.n101 VDD.t10 280.038
R49 VDD.n102 VDD.t20 280.038
R50 VDD.n108 VDD.t20 280.038
R51 VDD.n109 VDD.t6 280.038
R52 VDD.n115 VDD.t6 280.038
R53 VDD.n116 VDD.t0 280.038
R54 VDD.n122 VDD.t0 280.038
R55 VDD.n123 VDD.t22 280.038
R56 VDD.n129 VDD.t22 280.038
R57 VDD.n76 VDD.t14 280.038
R58 VDD.n75 VDD.t18 280.038
R59 VDD.n38 VDD.t18 280.038
R60 VDD.t2 VDD.n40 280.038
R61 VDD.n65 VDD.t2 280.038
R62 VDD.n64 VDD.t4 280.038
R63 VDD.n51 VDD.t4 280.038
R64 VDD.t12 VDD.n52 280.038
R65 VDD.n140 VDD.n4 255.526
R66 VDD.n96 VDD.n95 229.012
R67 VDD.n27 VDD.n26 229.012
R68 VDD.n55 VDD.n49 229.012
R69 VDD.n137 VDD.n136 184.957
R70 VDD.n52 VDD.n51 163.06
R71 VDD.n123 VDD.n122 161.287
R72 VDD.n102 VDD.n101 159.516
R73 VDD.n76 VDD.n75 159.516
R74 VDD.n116 VDD.n115 157.744
R75 VDD.n109 VDD.n108 155.97
R76 VDD.n40 VDD.n38 155.97
R77 VDD.n65 VDD.n64 155.97
R78 VDD.n125 VDD.n10 134.024
R79 VDD.n127 VDD.n10 134.024
R80 VDD.n126 VDD.n125 134.024
R81 VDD.n127 VDD.n126 134.024
R82 VDD.n118 VDD.n13 134.024
R83 VDD.n120 VDD.n13 134.024
R84 VDD.n119 VDD.n118 134.024
R85 VDD.n120 VDD.n119 134.024
R86 VDD.n111 VDD.n16 134.024
R87 VDD.n113 VDD.n16 134.024
R88 VDD.n112 VDD.n111 134.024
R89 VDD.n113 VDD.n112 134.024
R90 VDD.n104 VDD.n19 134.024
R91 VDD.n106 VDD.n19 134.024
R92 VDD.n105 VDD.n104 134.024
R93 VDD.n106 VDD.n105 134.024
R94 VDD.n99 VDD.n94 134.024
R95 VDD.n99 VDD.n98 134.024
R96 VDD.n98 VDD.n97 134.024
R97 VDD.n97 VDD.n94 134.024
R98 VDD.n24 VDD.n22 134.024
R99 VDD.n78 VDD.n24 134.024
R100 VDD.n79 VDD.n22 134.024
R101 VDD.n79 VDD.n78 134.024
R102 VDD.n73 VDD.n30 134.024
R103 VDD.n31 VDD.n30 134.024
R104 VDD.n73 VDD.n72 134.024
R105 VDD.n72 VDD.n31 134.024
R106 VDD.n35 VDD.n33 134.024
R107 VDD.n67 VDD.n35 134.024
R108 VDD.n68 VDD.n33 134.024
R109 VDD.n68 VDD.n67 134.024
R110 VDD.n62 VDD.n43 134.024
R111 VDD.n44 VDD.n43 134.024
R112 VDD.n62 VDD.n61 134.024
R113 VDD.n61 VDD.n44 134.024
R114 VDD.n53 VDD.n46 134.024
R115 VDD.n57 VDD.n46 134.024
R116 VDD.n53 VDD.n47 134.024
R117 VDD.n57 VDD.n47 134.024
R118 VDD.n132 VDD.n7 118.213
R119 VDD.n134 VDD.n7 118.213
R120 VDD.n133 VDD.n132 118.213
R121 VDD.n134 VDD.n133 118.213
R122 VDD.n142 VDD.n1 118.213
R123 VDD.n142 VDD.n2 118.213
R124 VDD.n138 VDD.n1 118.213
R125 VDD.n138 VDD.n2 118.213
R126 VDD.n144 VDD.t17 68.3354
R127 VDD.n82 VDD.t9 68.3354
R128 VDD.n81 VDD.t15 34.3985
R129 VDD.n32 VDD.t19 34.3985
R130 VDD.n70 VDD.t3 34.3985
R131 VDD.n45 VDD.t5 34.3985
R132 VDD.n59 VDD.t13 34.3985
R133 VDD.n84 VDD.t23 34.3985
R134 VDD.n86 VDD.t1 34.3985
R135 VDD.n88 VDD.t7 34.3985
R136 VDD.n90 VDD.t21 34.3985
R137 VDD.n92 VDD.t11 34.3985
R138 VDD.n93 VDD.n81 3.74141
R139 VDD.n143 VDD.n0 0.515806
R140 VDD.n80 VDD 0.26425
R141 VDD.n71 VDD 0.26425
R142 VDD.n69 VDD 0.26425
R143 VDD.n60 VDD 0.26425
R144 VDD.n58 VDD 0.26425
R145 VDD VDD.n85 0.2455
R146 VDD VDD.n91 0.24425
R147 VDD VDD.n87 0.243
R148 VDD VDD.n89 0.24175
R149 VDD.n92 VDD 0.20675
R150 VDD.n90 VDD 0.20675
R151 VDD.n88 VDD 0.20675
R152 VDD.n86 VDD 0.20675
R153 VDD VDD.n144 0.203306
R154 VDD VDD.n82 0.200755
R155 VDD.n84 VDD.n83 0.19425
R156 VDD VDD.n59 0.18925
R157 VDD.n32 VDD 0.18675
R158 VDD VDD.n70 0.18425
R159 VDD.n45 VDD 0.18425
R160 VDD.n81 VDD.n80 0.058
R161 VDD.n71 VDD.n32 0.058
R162 VDD.n70 VDD.n69 0.058
R163 VDD.n60 VDD.n45 0.058
R164 VDD.n59 VDD.n58 0.058
R165 VDD.n93 VDD.n92 0.058
R166 VDD.n91 VDD.n90 0.058
R167 VDD.n89 VDD.n88 0.058
R168 VDD.n87 VDD.n86 0.058
R169 VDD.n85 VDD.n84 0.058
R170 VDD.n82 VDD.n0 0.0566224
R171 VDD.n144 VDD.n143 0.0566224
R172 VDD.n139 VDD.n138 0.0349892
R173 VDD.n133 VDD.n6 0.0349892
R174 VDD.n6 VDD.t8 0.0349892
R175 VDD.n105 VDD.n18 0.0349892
R176 VDD.n18 VDD.t20 0.0349892
R177 VDD.n112 VDD.n15 0.0349892
R178 VDD.n15 VDD.t6 0.0349892
R179 VDD.n119 VDD.n12 0.0349892
R180 VDD.n12 VDD.t0 0.0349892
R181 VDD.n126 VDD.n9 0.0349892
R182 VDD.n9 VDD.t22 0.0349892
R183 VDD.n98 VDD.n21 0.0349892
R184 VDD.n21 VDD.t10 0.0349892
R185 VDD.n43 VDD.n41 0.0349892
R186 VDD.n41 VDD.t4 0.0349892
R187 VDD.n36 VDD.n35 0.0349892
R188 VDD.t2 VDD.n36 0.0349892
R189 VDD.n30 VDD.n28 0.0349892
R190 VDD.n28 VDD.t18 0.0349892
R191 VDD.n25 VDD.n24 0.0349892
R192 VDD.t14 VDD.n25 0.0349892
R193 VDD.n54 VDD.n53 0.0349892
R194 VDD.t12 VDD.n54 0.0349892
R195 VDD.n4 VDD.n2 0.0286326
R196 VDD.n3 VDD.n1 0.0286326
R197 VDD.n137 VDD.n3 0.0286326
R198 VDD.n135 VDD.n134 0.0286326
R199 VDD.n136 VDD.n135 0.0286326
R200 VDD.n132 VDD.n131 0.0286326
R201 VDD.n131 VDD.n130 0.0286326
R202 VDD.n140 VDD.n139 0.0275362
R203 VDD.n107 VDD.n106 0.018623
R204 VDD.n108 VDD.n107 0.018623
R205 VDD.n104 VDD.n103 0.018623
R206 VDD.n103 VDD.n102 0.018623
R207 VDD.n114 VDD.n113 0.018623
R208 VDD.n115 VDD.n114 0.018623
R209 VDD.n111 VDD.n110 0.018623
R210 VDD.n110 VDD.n109 0.018623
R211 VDD.n121 VDD.n120 0.018623
R212 VDD.n122 VDD.n121 0.018623
R213 VDD.n118 VDD.n117 0.018623
R214 VDD.n117 VDD.n116 0.018623
R215 VDD.n128 VDD.n127 0.018623
R216 VDD.n129 VDD.n128 0.018623
R217 VDD.n125 VDD.n124 0.018623
R218 VDD.n124 VDD.n123 0.018623
R219 VDD.n100 VDD.n99 0.018623
R220 VDD.n101 VDD.n100 0.018623
R221 VDD.n97 VDD.n96 0.018623
R222 VDD.n50 VDD.n44 0.018623
R223 VDD.n51 VDD.n50 0.018623
R224 VDD.n63 VDD.n62 0.018623
R225 VDD.n64 VDD.n63 0.018623
R226 VDD.n67 VDD.n66 0.018623
R227 VDD.n66 VDD.n65 0.018623
R228 VDD.n39 VDD.n33 0.018623
R229 VDD.n40 VDD.n39 0.018623
R230 VDD.n37 VDD.n31 0.018623
R231 VDD.n38 VDD.n37 0.018623
R232 VDD.n74 VDD.n73 0.018623
R233 VDD.n75 VDD.n74 0.018623
R234 VDD.n78 VDD.n77 0.018623
R235 VDD.n77 VDD.n76 0.018623
R236 VDD.n26 VDD.n22 0.018623
R237 VDD.n48 VDD.n46 0.018623
R238 VDD.n52 VDD.n48 0.018623
R239 VDD.n49 VDD.n47 0.018623
R240 VDD.n83 VDD 0.013005
R241 VDD.n83 VDD 0.013
R242 VDD.t16 VDD.n140 0.00895217
R243 VDD.n42 VDD.t4 0.00380159
R244 VDD.t2 VDD.n34 0.00380159
R245 VDD.n29 VDD.t18 0.00380159
R246 VDD.n57 VDD.n56 0.00380159
R247 VDD.n61 VDD.n42 0.00380159
R248 VDD.n68 VDD.n34 0.00380159
R249 VDD.n72 VDD.n29 0.00380159
R250 VDD.n79 VDD.n23 0.00380159
R251 VDD.n94 VDD.n20 0.00380159
R252 VDD.n19 VDD.n17 0.00380159
R253 VDD.n17 VDD.t20 0.00380159
R254 VDD.n16 VDD.n14 0.00380159
R255 VDD.n14 VDD.t6 0.00380159
R256 VDD.n13 VDD.n11 0.00380159
R257 VDD.n11 VDD.t0 0.00380159
R258 VDD.n10 VDD.n8 0.00380159
R259 VDD.n8 VDD.t22 0.00380159
R260 VDD.n7 VDD.n5 0.00380159
R261 VDD.n5 VDD.t8 0.00380159
R262 VDD.n142 VDD.n141 0.00380159
R263 VDD.n141 VDD.t16 0.00380159
R264 VDD.n95 VDD.n20 0.00369982
R265 VDD.n27 VDD.n23 0.00369982
R266 VDD.n56 VDD.n55 0.00369982
R267 VDD.n58 VDD.n57 0.00233287
R268 VDD.n61 VDD.n60 0.00233287
R269 VDD.n69 VDD.n68 0.00233287
R270 VDD.n72 VDD.n71 0.00233287
R271 VDD.n80 VDD.n79 0.00233287
R272 VDD.n94 VDD.n93 0.00233287
R273 VDD.n91 VDD.n19 0.00233287
R274 VDD.n89 VDD.n16 0.00233287
R275 VDD.n87 VDD.n13 0.00233287
R276 VDD.n85 VDD.n10 0.00233287
R277 VDD.n7 VDD.n0 0.00233287
R278 VDD.n143 VDD.n142 0.00233287
R279 VDD.t14 VDD.n27 0.00160176
R280 VDD.n55 VDD.t12 0.00160176
R281 VDD.n95 VDD.t10 0.00160176
R282 CLK.n1 CLK.t2 155.125
R283 CLK.n2 CLK.t3 140.486
R284 CLK.n0 CLK.t0 42.4671
R285 CLK.n0 CLK.t1 35.198
R286 CLK CLK.n2 4.52884
R287 CLK.n2 CLK.n1 0.388431
R288 CLK CLK.n0 0.340778
R289 CLK.n1 CLK 0.274538
R290 VSS.n97 VSS.n96 451.92
R291 VSS.n52 VSS.n51 446.954
R292 VSS.n62 VSS.n61 437.021
R293 VSS.n83 VSS.n82 437.021
R294 VSS.n128 VSS.n121 116.329
R295 VSS.n128 VSS.n127 116.329
R296 VSS.n104 VSS.n99 116.329
R297 VSS.n104 VSS.n103 116.329
R298 VSS.n94 VSS.n15 116.329
R299 VSS.n93 VSS.n18 116.329
R300 VSS.n94 VSS.n93 116.329
R301 VSS.n59 VSS.n22 116.329
R302 VSS.n72 VSS.n22 116.329
R303 VSS.n72 VSS.n71 116.329
R304 VSS.n29 VSS.n27 116.329
R305 VSS.n64 VSS.n29 116.329
R306 VSS.n65 VSS.n64 116.329
R307 VSS.n35 VSS.n33 116.329
R308 VSS.n40 VSS.n35 116.329
R309 VSS.n40 VSS.n39 116.329
R310 VSS.n49 VSS.n43 116.329
R311 VSS.n48 VSS.n46 116.329
R312 VSS.n49 VSS.n48 116.329
R313 VSS.n57 VSS.n31 116.329
R314 VSS.n56 VSS.n54 116.329
R315 VSS.n57 VSS.n56 116.329
R316 VSS.n77 VSS.n75 116.329
R317 VSS.n80 VSS.n77 116.329
R318 VSS.n80 VSS.n79 116.329
R319 VSS.n89 VSS.n85 116.329
R320 VSS.n117 VSS.n110 116.329
R321 VSS.n117 VSS.n112 116.329
R322 VSS.n10 VSS.n4 116.329
R323 VSS.n10 VSS.n2 116.329
R324 VSS.n38 VSS.t12 41.7657
R325 VSS.n107 VSS.t14 41.7387
R326 VSS.n37 VSS.t9 41.7354
R327 VSS.n67 VSS.t17 41.7354
R328 VSS.n69 VSS.t7 41.7354
R329 VSS.n91 VSS.t1 41.7354
R330 VSS.n106 VSS.t18 41.7354
R331 VSS.n0 VSS.t11 41.7354
R332 VSS.n20 VSS.t6 41.7354
R333 VSS.n68 VSS.t3 41.7354
R334 VSS.n24 VSS.t16 41.7354
R335 VSS.n96 VSS.n13 4.96664
R336 VSS.n129 VSS.n118 0.515806
R337 VSS VSS.n129 0.254327
R338 VSS.n107 VSS 0.198204
R339 VSS.n87 VSS.n86 0.10956
R340 VSS.t5 VSS.n87 0.10956
R341 VSS.n79 VSS.n78 0.10956
R342 VSS.n56 VSS.n55 0.10956
R343 VSS.n48 VSS.n47 0.10956
R344 VSS.n35 VSS.n34 0.10956
R345 VSS.n29 VSS.n28 0.10956
R346 VSS.n22 VSS.n21 0.10956
R347 VSS.n15 VSS.n14 0.10956
R348 VSS.n8 VSS.n7 0.10956
R349 VSS.t10 VSS.n8 0.10956
R350 VSS.n123 VSS.n122 0.10956
R351 VSS.t4 VSS.n123 0.10956
R352 VSS.n114 VSS.n113 0.10956
R353 VSS.n6 VSS.n5 0.10956
R354 VSS.t10 VSS.n6 0.10956
R355 VSS.n37 VSS 0.106814
R356 VSS VSS.n67 0.106814
R357 VSS.n69 VSS 0.106814
R358 VSS VSS.n106 0.106814
R359 VSS.n91 VSS 0.10617
R360 VSS VSS.n0 0.0958608
R361 VSS VSS.n24 0.0952165
R362 VSS.n112 VSS.n111 0.0944005
R363 VSS.n12 VSS.n11 0.0944005
R364 VSS.n13 VSS.n12 0.0944005
R365 VSS.n85 VSS.n84 0.0944005
R366 VSS.n84 VSS.n83 0.0944005
R367 VSS.n81 VSS.n80 0.0944005
R368 VSS.n82 VSS.n81 0.0944005
R369 VSS.n75 VSS.n74 0.0944005
R370 VSS.n58 VSS.n57 0.0944005
R371 VSS.n62 VSS.n58 0.0944005
R372 VSS.n54 VSS.n53 0.0944005
R373 VSS.n53 VSS.n52 0.0944005
R374 VSS.n50 VSS.n49 0.0944005
R375 VSS.n51 VSS.n50 0.0944005
R376 VSS.n46 VSS.n45 0.0944005
R377 VSS.n45 VSS.n44 0.0944005
R378 VSS.n41 VSS.n40 0.0944005
R379 VSS.n51 VSS.n41 0.0944005
R380 VSS.n33 VSS.n32 0.0944005
R381 VSS.n64 VSS.n63 0.0944005
R382 VSS.n63 VSS.n62 0.0944005
R383 VSS.n27 VSS.n26 0.0944005
R384 VSS.n73 VSS.n72 0.0944005
R385 VSS.n82 VSS.n73 0.0944005
R386 VSS.n60 VSS.n59 0.0944005
R387 VSS.n61 VSS.n60 0.0944005
R388 VSS.n95 VSS.n94 0.0944005
R389 VSS.n96 VSS.n95 0.0944005
R390 VSS.n18 VSS.n17 0.0944005
R391 VSS.n17 VSS.n16 0.0944005
R392 VSS.n103 VSS.n102 0.0944005
R393 VSS.n102 VSS.n101 0.0944005
R394 VSS.n99 VSS.n98 0.0944005
R395 VSS.n98 VSS.n97 0.0944005
R396 VSS.n127 VSS.n126 0.0944005
R397 VSS.n126 VSS.n125 0.0944005
R398 VSS.n121 VSS.n120 0.0944005
R399 VSS.n120 VSS.n119 0.0944005
R400 VSS.n110 VSS.n109 0.0944005
R401 VSS.n109 VSS.n108 0.0944005
R402 VSS.n4 VSS.n3 0.0944005
R403 VSS.n2 VSS.n1 0.0944005
R404 VSS.n68 VSS 0.0939278
R405 VSS VSS.n20 0.0939278
R406 VSS.n115 VSS.n114 0.0768221
R407 VSS.n118 VSS.n107 0.0591735
R408 VSS.t13 VSS.n115 0.0342337
R409 VSS.n38 VSS.n37 0.0307835
R410 VSS.n66 VSS.n24 0.0307835
R411 VSS.n67 VSS.n66 0.0307835
R412 VSS.n70 VSS.n68 0.0307835
R413 VSS.n70 VSS.n69 0.0307835
R414 VSS.n90 VSS.n20 0.0307835
R415 VSS.n92 VSS.n91 0.0307835
R416 VSS.n105 VSS.n0 0.0307835
R417 VSS.n106 VSS.n105 0.0307835
R418 VSS.n36 VSS.t8 0.0039133
R419 VSS.n25 VSS.t15 0.0039133
R420 VSS.n23 VSS.t2 0.0039133
R421 VSS.n19 VSS.t0 0.0039133
R422 VSS.n124 VSS.t4 0.0039133
R423 VSS.n116 VSS.t13 0.0039133
R424 VSS.n9 VSS.t10 0.0039133
R425 VSS.n10 VSS.n9 0.0039133
R426 VSS.n89 VSS.n88 0.0039133
R427 VSS.n88 VSS.t5 0.0039133
R428 VSS.n77 VSS.n76 0.0039133
R429 VSS.n31 VSS.n30 0.0039133
R430 VSS.n43 VSS.n42 0.0039133
R431 VSS.n39 VSS.n36 0.0039133
R432 VSS.n65 VSS.n25 0.0039133
R433 VSS.n71 VSS.n23 0.0039133
R434 VSS.n93 VSS.n19 0.0039133
R435 VSS.n104 VSS.n100 0.0039133
R436 VSS.n128 VSS.n124 0.0039133
R437 VSS.n117 VSS.n116 0.0039133
R438 VSS.n105 VSS.n10 0.00233287
R439 VSS.n90 VSS.n89 0.00233287
R440 VSS.n39 VSS.n38 0.00233287
R441 VSS.n66 VSS.n65 0.00233287
R442 VSS.n71 VSS.n70 0.00233287
R443 VSS.n93 VSS.n92 0.00233287
R444 VSS.n105 VSS.n104 0.00233287
R445 VSS.n129 VSS.n128 0.00233287
R446 VSS.n118 VSS.n117 0.00233287
R447 VSS.n92 VSS.n90 0.00114433
R448 EN_CLK.n0 EN_CLK.t0 155.132
R449 EN_CLK.n0 EN_CLK.t1 140.864
R450 EN_CLK EN_CLK.n0 0.382411
C0 x2.Vin x4.Vin 3.23e-19
C1 x9.Vin x5.Vin 9.41e-20
C2 x9.Vin x4.Vin 0.0031f
C3 x5.Vin x6.Vin 0.184f
C4 a_1692_1940# CLK 0.0379f
C5 x3.Vin CLK 0.0052f
C6 x2.Vin x11.Vin 0.0031f
C7 x2.Vin x6.Vin 2.59e-20
C8 x9.Vout x4.Vin 9.79e-20
C9 VDD a_1692_1940# 0.00823f
C10 x3.Vin VDD 0.634f
C11 VDD CLK 0.63f
C12 x6.Vin x7.Vin 0.177f
C13 EN_CLK a_1692_1940# 0.0121f
C14 EN_CLK CLK 0.0282f
C15 x9.Vout x11.Vin 0.184f
C16 EN_CLK VDD 0.268f
C17 x9.Vout x9.Vin 0.184f
C18 x8.Vin CLK 8.11e-20
C19 VDD x8.Vin 0.637f
C20 x4.Vin x3.Vin 0.184f
C21 x5.Vin CLK 2.68e-19
C22 x4.Vin CLK 6.64e-19
C23 x5.Vin VDD 0.633f
C24 x4.Vin VDD 0.633f
C25 x2.Vin a_1692_1940# 0.108f
C26 x2.Vin x3.Vin 0.181f
C27 x2.Vin CLK 0.411f
C28 x3.Vin x11.Vin 9.79e-20
C29 x2.Vin VDD 0.798f
C30 CLK x11.Vin 0.177f
C31 x9.Vin CLK 4.98e-19
C32 VDD x7.Vin 1.18f
C33 x2.Vin EN_CLK 0.0822f
C34 VDD x11.Vin 0.628f
C35 x9.Vin VDD 0.633f
C36 x5.Vin x8.Vin 0.0031f
C37 VDD x6.Vin 0.63f
C38 x9.Vout x3.Vin 0.0031f
C39 x9.Vout CLK 0.00102f
C40 x9.Vout VDD 0.633f
C41 x4.Vin x5.Vin 0.184f
C42 x8.Vin x7.Vin 0.18f
C43 x9.Vin x8.Vin 0.184f
C44 x8.Vin x6.Vin 9.41e-20
C45 x2.Vin x5.Vin 1.46e-19
C46 x8.Vin 0 0.583f
C47 x9.Vin 0 0.582f
C48 x9.Vout 0 0.582f
C49 x11.Vin 0 0.598f
C50 a_1692_1940# 0 0.372f
C51 x7.Vin 0 0.853f
C52 x6.Vin 0 0.597f
C53 x5.Vin 0 0.582f
C54 x4.Vin 0 0.582f
C55 x3.Vin 0 0.583f
C56 CLK 0 1.14f
C57 x2.Vin 0 0.719f
C58 EN_CLK 0 0.413f
C59 VDD 0 12.1f
.ends

