magic
tech sky130A
magscale 1 2
timestamp 1691650988
<< nwell >>
rect 478 396 1304 848
<< pwell >>
rect 482 -204 1308 238
<< nmos >>
rect 678 -56 708 28
rect 1082 -56 1112 28
<< pmos >>
rect 674 616 704 700
rect 1078 616 1108 700
<< ndiff >>
rect 620 16 678 28
rect 620 -44 632 16
rect 666 -44 678 16
rect 620 -56 678 -44
rect 708 16 766 28
rect 708 -44 720 16
rect 754 -44 766 16
rect 708 -56 766 -44
rect 1024 16 1082 28
rect 1024 -44 1036 16
rect 1070 -44 1082 16
rect 1024 -56 1082 -44
rect 1112 16 1170 28
rect 1112 -44 1124 16
rect 1158 -44 1170 16
rect 1112 -56 1170 -44
<< pdiff >>
rect 616 688 674 700
rect 616 628 628 688
rect 662 628 674 688
rect 616 616 674 628
rect 704 688 762 700
rect 704 628 716 688
rect 750 628 762 688
rect 704 616 762 628
rect 1020 688 1078 700
rect 1020 628 1032 688
rect 1066 628 1078 688
rect 1020 616 1078 628
rect 1108 688 1166 700
rect 1108 628 1120 688
rect 1154 628 1166 688
rect 1108 616 1166 628
<< ndiffc >>
rect 632 -44 666 16
rect 720 -44 754 16
rect 1036 -44 1070 16
rect 1124 -44 1158 16
<< pdiffc >>
rect 628 628 662 688
rect 716 628 750 688
rect 1032 628 1066 688
rect 1120 628 1154 688
<< psubdiff >>
rect 518 168 614 202
rect 772 168 868 202
rect 518 106 552 168
rect 834 106 868 168
rect 518 -134 552 -72
rect 834 -134 868 -72
rect 518 -168 614 -134
rect 772 -168 868 -134
rect 922 168 1018 202
rect 1176 168 1272 202
rect 922 106 956 168
rect 1238 106 1272 168
rect 922 -134 956 -72
rect 1238 -134 1272 -72
rect 922 -168 1018 -134
rect 1176 -168 1272 -134
<< nsubdiff >>
rect 514 778 610 812
rect 768 778 864 812
rect 514 715 548 778
rect 830 715 864 778
rect 514 466 548 529
rect 830 466 864 529
rect 514 432 610 466
rect 768 432 864 466
rect 918 778 1014 812
rect 1172 778 1268 812
rect 918 715 952 778
rect 1234 715 1268 778
rect 918 466 952 529
rect 1234 466 1268 529
rect 918 432 1014 466
rect 1172 432 1268 466
<< psubdiffcont >>
rect 614 168 772 202
rect 518 -72 552 106
rect 834 -72 868 106
rect 614 -168 772 -134
rect 1018 168 1176 202
rect 922 -72 956 106
rect 1238 -72 1272 106
rect 1018 -168 1176 -134
<< nsubdiffcont >>
rect 610 778 768 812
rect 514 529 548 715
rect 830 529 864 715
rect 610 432 768 466
rect 1014 778 1172 812
rect 918 529 952 715
rect 1234 529 1268 715
rect 1014 432 1172 466
<< poly >>
rect 674 700 704 726
rect 674 585 704 616
rect 656 569 722 585
rect 656 535 672 569
rect 706 535 722 569
rect 656 519 722 535
rect 1078 700 1108 726
rect 1078 585 1108 616
rect 1060 569 1126 585
rect 1060 535 1076 569
rect 1110 535 1126 569
rect 1060 519 1126 535
rect 660 100 726 116
rect 660 66 676 100
rect 710 66 726 100
rect 660 50 726 66
rect 678 28 708 50
rect 678 -82 708 -56
rect 1064 100 1130 116
rect 1064 66 1080 100
rect 1114 66 1130 100
rect 1064 50 1130 66
rect 1082 28 1112 50
rect 1082 -82 1112 -56
<< polycont >>
rect 672 535 706 569
rect 1076 535 1110 569
rect 676 66 710 100
rect 1080 66 1114 100
<< locali >>
rect 514 778 610 812
rect 768 778 864 812
rect 514 715 548 778
rect 830 715 864 778
rect 628 688 662 704
rect 628 612 662 628
rect 716 688 750 704
rect 716 612 750 628
rect 656 535 672 569
rect 706 535 722 569
rect 514 466 548 529
rect 830 466 864 529
rect 514 432 610 466
rect 768 432 864 466
rect 918 778 1014 812
rect 1172 778 1268 812
rect 918 715 952 778
rect 1234 715 1268 778
rect 1032 688 1066 704
rect 1032 612 1066 628
rect 1120 688 1154 704
rect 1120 612 1154 628
rect 1060 535 1076 569
rect 1110 535 1126 569
rect 918 466 952 529
rect 1234 466 1268 529
rect 918 432 1014 466
rect 1172 432 1268 466
rect 518 168 614 202
rect 772 168 868 202
rect 518 106 552 168
rect 834 106 868 168
rect 660 66 676 100
rect 710 66 726 100
rect 632 16 666 32
rect 632 -60 666 -44
rect 720 16 754 32
rect 720 -60 754 -44
rect 518 -134 552 -72
rect 834 -134 868 -72
rect 518 -168 614 -134
rect 772 -168 868 -134
rect 922 168 1018 202
rect 1176 168 1272 202
rect 922 106 956 168
rect 1238 106 1272 168
rect 1064 66 1080 100
rect 1114 66 1130 100
rect 1036 16 1070 32
rect 1036 -60 1070 -44
rect 1124 16 1158 32
rect 1124 -60 1158 -44
rect 922 -134 956 -72
rect 1238 -134 1272 -72
rect 922 -168 1018 -134
rect 1176 -168 1272 -134
<< viali >>
rect 610 778 768 812
rect 628 628 662 688
rect 716 628 750 688
rect 672 535 706 569
rect 1014 778 1172 812
rect 1032 628 1066 688
rect 1120 628 1154 688
rect 1076 535 1110 569
rect 676 66 710 100
rect 632 -44 666 16
rect 720 -44 754 16
rect 614 -168 772 -134
rect 1080 66 1114 100
rect 1036 -44 1070 16
rect 1124 -44 1158 16
rect 1018 -168 1176 -134
<< metal1 >>
rect 478 812 1304 848
rect 478 778 610 812
rect 768 778 1014 812
rect 1172 778 1304 812
rect 478 750 1304 778
rect 628 700 662 750
rect 1120 700 1154 750
rect 622 688 668 700
rect 622 628 628 688
rect 662 628 668 688
rect 622 616 668 628
rect 710 688 756 700
rect 710 628 716 688
rect 750 662 756 688
rect 1026 688 1072 700
rect 1026 662 1032 688
rect 750 628 1032 662
rect 1066 628 1072 688
rect 710 622 1072 628
rect 710 616 756 622
rect 670 575 716 576
rect 660 569 718 575
rect 660 535 672 569
rect 706 535 718 569
rect 660 529 718 535
rect 670 106 716 529
rect 868 372 914 622
rect 1026 616 1072 622
rect 1114 688 1160 700
rect 1114 628 1120 688
rect 1154 628 1160 688
rect 1114 616 1160 628
rect 1064 569 1122 575
rect 1064 535 1076 569
rect 1110 535 1122 569
rect 1064 529 1122 535
rect 854 366 930 372
rect 854 302 860 366
rect 924 302 930 366
rect 854 296 930 302
rect 1070 106 1116 529
rect 1176 360 1240 366
rect 1176 308 1182 360
rect 1234 308 1240 360
rect 1176 302 1240 308
rect 664 100 722 106
rect 664 66 676 100
rect 710 66 722 100
rect 664 60 722 66
rect 1068 100 1126 106
rect 1068 66 1080 100
rect 1114 66 1126 100
rect 1068 60 1126 66
rect 1070 58 1116 60
rect 1192 28 1228 302
rect 626 16 672 28
rect 626 -44 632 16
rect 666 -44 672 16
rect 626 -56 672 -44
rect 714 16 760 28
rect 714 -44 720 16
rect 754 6 760 16
rect 1030 16 1076 28
rect 1030 6 1036 16
rect 754 -34 1036 6
rect 754 -44 760 -34
rect 714 -56 760 -44
rect 1030 -44 1036 -34
rect 1070 -44 1076 16
rect 1030 -56 1076 -44
rect 1118 16 1228 28
rect 1118 -44 1124 16
rect 1158 -12 1228 16
rect 1158 -44 1164 -12
rect 1118 -56 1164 -44
rect 628 -108 666 -56
rect 482 -134 1308 -108
rect 482 -168 614 -134
rect 772 -168 1018 -134
rect 1176 -168 1308 -134
rect 482 -206 1308 -168
<< via1 >>
rect 860 302 924 366
rect 1182 308 1234 360
<< metal2 >>
rect 854 366 930 372
rect 854 302 860 366
rect 924 356 930 366
rect 1176 360 1240 366
rect 1176 356 1182 360
rect 924 314 1182 356
rect 924 302 930 314
rect 1176 308 1182 314
rect 1234 356 1240 360
rect 1234 314 1312 356
rect 1234 308 1240 314
rect 1176 302 1240 308
rect 854 296 930 302
<< labels >>
flabel space 670 60 716 576 0 FreeSans 160 0 0 0 A
port 0 nsew
flabel space 1070 58 1116 575 0 FreeSans 160 0 0 0 B
port 1 nsew
flabel metal2 1234 314 1312 356 0 FreeSans 160 0 0 0 OUT
port 2 nsew
flabel metal1 478 812 1304 848 0 FreeSans 160 0 0 0 VDD
port 3 nsew
flabel metal1 482 -206 1308 -168 0 FreeSans 160 0 0 0 VSS
port 5 nsew
<< end >>
