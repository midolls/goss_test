magic
tech sky130A
magscale 1 2
timestamp 1691735525
<< metal1 >>
rect 4304 2762 4504 2766
rect 1474 2696 1580 2760
rect 4304 2678 4524 2762
rect 1464 2288 1570 2352
rect 2202 2216 2314 2250
rect 4322 2248 4358 2250
rect 4322 2214 4394 2248
rect 2052 2172 2116 2178
rect 2052 2120 2058 2172
rect 2110 2120 2116 2172
rect 2052 2114 2116 2120
rect 1474 1806 1582 1870
rect 2048 1378 2112 1384
rect 2048 1326 2054 1378
rect 2108 1368 2112 1378
rect 4354 1368 4394 2214
rect 2108 1332 2280 1368
rect 4322 1334 4394 1368
rect 4322 1332 4358 1334
rect 2108 1326 2112 1332
rect 2048 1320 2112 1326
rect 4426 904 4524 2678
rect 4304 816 4524 904
<< via1 >>
rect 2058 2120 2110 2172
rect 2054 1326 2108 1378
<< metal2 >>
rect 2052 2172 2116 2178
rect 2052 2120 2058 2172
rect 2110 2120 2116 2172
rect 2052 2114 2116 2120
rect 2058 1384 2106 2114
rect 2048 1378 2112 1384
rect 2048 1326 2054 1378
rect 2108 1326 2112 1378
rect 2048 1320 2112 1326
use nand  x1
timestamp 1691733244
transform 1 0 988 0 1 1924
box 478 -134 1312 848
use inverter  x2
timestamp 1691733642
transform 1 0 1966 0 1 1800
box 314 -10 738 970
use inverter  x3
timestamp 1691733642
transform 1 0 2373 0 1 1800
box 314 -10 738 970
use inverter  x4
timestamp 1691733642
transform 1 0 2778 0 1 1800
box 314 -10 738 970
use inverter  x5
timestamp 1691733642
transform 1 0 3182 0 1 1800
box 314 -10 738 970
use inverter  x6
timestamp 1691733642
transform 1 0 3588 0 1 1800
box 314 -10 738 970
use inverter  x7
timestamp 1691733642
transform -1 0 4640 0 -1 1782
box 314 -10 738 970
use inverter  x8
timestamp 1691733642
transform -1 0 4234 0 -1 1782
box 314 -10 738 970
use inverter  x9
timestamp 1691733642
transform -1 0 3830 0 -1 1782
box 314 -10 738 970
use inverter  x10
timestamp 1691733642
transform -1 0 3426 0 -1 1782
box 314 -10 738 970
use inverter  x11
timestamp 1691733642
transform -1 0 3018 0 -1 1782
box 314 -10 738 970
<< labels >>
flabel metal1 2154 1332 2250 1362 0 FreeSans 160 0 0 0 CLK
port 5 nsew
flabel metal1 1474 2696 1580 2760 0 FreeSans 160 0 0 0 VDD
port 0 nsew
flabel metal1 1476 1806 1582 1870 0 FreeSans 160 0 0 0 VSS
port 1 nsew
flabel metal1 1464 2288 1570 2352 0 FreeSans 160 0 0 0 EN_CLK
port 7 nsew
<< end >>
