* NGSPICE file created from inverter_flat.ext - technology: sky130A

.subckt inverter_flat Vin Vout VDD VSS
X0 Vout.t1 Vin.t0 VSS.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1 Vout.t0 Vin.t1 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
R0 Vin.n0 Vin.t1 222.611
R1 Vin Vin.t0 140.625
R2 Vin.n0 Vin 0.6255
R3 Vin Vin.n0 0.038
R4 VSS.n8 VSS.n7 90.2269
R5 VSS.n14 VSS.n13 81.0463
R6 VSS.n11 VSS.t1 41.7354
R7 VSS.n15 VSS.n14 9.3005
R8 VSS VSS.n15 0.152286
R9 VSS.n1 VSS.n0 0.10956
R10 VSS.n13 VSS.n12 0.0944005
R11 VSS.n7 VSS.n6 0.0944005
R12 VSS.n2 VSS.n1 0.0592926
R13 VSS.n15 VSS.n11 0.0591735
R14 VSS.n11 VSS.n10 0.0553469
R15 VSS.t0 VSS.n2 0.0520137
R16 VSS.n10 VSS.n8 0.00690386
R17 VSS.n5 VSS.n4 0.0039133
R18 VSS.n8 VSS.n5 0.00366545
R19 VSS.n4 VSS.n3 0.00282082
R20 VSS.n3 VSS.t0 0.00259248
R21 VSS.n10 VSS.n9 0.000572701
R22 Vout Vout.t1 42.4673
R23 Vout Vout.t0 35.2375
R24 VDD.n8 VDD.n1 106.049
R25 VDD.n12 VDD.n11 98.7195
R26 VDD.n9 VDD.t1 34.3985
R27 VDD.n13 VDD.n12 9.3005
R28 VDD VDD.n13 0.148
R29 VDD.n13 VDD.n9 0.05925
R30 VDD.n9 VDD.n8 0.0588938
R31 VDD.n3 VDD.n2 0.0349892
R32 VDD.t0 VDD.n3 0.0349892
R33 VDD.n11 VDD.n10 0.018623
R34 VDD.n1 VDD.n0 0.018623
R35 VDD.t0 VDD.n4 0.0135718
R36 VDD.n6 VDD.n5 0.00383554
R37 VDD.n7 VDD.n6 0.00380159
R38 VDD.n5 VDD.t0 0.00163201
R39 VDD.n8 VDD.n7 0.00142302
C0 VDD Vin 0.25f
C1 VDD Vout 0.326f
C2 Vout Vin 0.166f
.ends

