* NGSPICE file created from nand.ext - technology: sky130A

.subckt nand OUT A B VDD VSS
X0 VDD.t3 B.t0 OUT.t2 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1 OUT.t1 B.t1 a_704_16# VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X2 OUT.t0 A.t0 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X3 a_704_16# A.t1 VSS.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
R0 B.n0 B.t0 155.125
R1 B.n0 B.t1 140.874
R2 B B.n0 0.274538
R3 OUT.n0 OUT.t2 68.4216
R4 OUT.n0 OUT.t0 68.4216
R5 OUT.n1 OUT.t1 44.425
R6 OUT.n1 OUT.n0 1.71365
R7 OUT OUT.n1 0.0512812
R8 VDD.n20 VDD.n13 118.213
R9 VDD.n20 VDD.n15 118.213
R10 VDD.n9 VDD.n4 118.213
R11 VDD.n9 VDD.n1 118.213
R12 VDD.n10 VDD.t3 68.3915
R13 VDD.n22 VDD.t1 68.3354
R14 VDD.n21 VDD.n10 0.515806
R15 VDD VDD.n22 0.21351
R16 VDD.n22 VDD.n21 0.0566224
R17 VDD.n17 VDD.n16 0.0349892
R18 VDD.n6 VDD.n5 0.0349892
R19 VDD.t2 VDD.n6 0.0349892
R20 VDD.n15 VDD.n14 0.0286326
R21 VDD.n13 VDD.n12 0.0286326
R22 VDD.n12 VDD.n11 0.0286326
R23 VDD.n4 VDD.n3 0.0286326
R24 VDD.n3 VDD.n2 0.0286326
R25 VDD.n1 VDD.n0 0.0286326
R26 VDD.n18 VDD.n17 0.0275362
R27 VDD.t0 VDD.n18 0.00895217
R28 VDD.n9 VDD.n8 0.00380159
R29 VDD.n20 VDD.n19 0.00380159
R30 VDD.n19 VDD.t0 0.00380159
R31 VDD.n8 VDD.n7 0.00354032
R32 VDD.n10 VDD.n9 0.00233287
R33 VDD.n21 VDD.n20 0.00233287
R34 VDD.n7 VDD.t2 0.00176126
R35 VSS.n19 VSS.n12 116.329
R36 VSS.n19 VSS.n14 116.329
R37 VSS.n9 VSS.n1 116.329
R38 VSS.n9 VSS.n4 116.329
R39 VSS.n21 VSS.t1 41.7387
R40 VSS.n20 VSS.n9 0.517639
R41 VSS VSS.n21 0.210959
R42 VSS.n16 VSS.n15 0.10956
R43 VSS.n6 VSS.n5 0.10956
R44 VSS.n14 VSS.n13 0.0944005
R45 VSS.n12 VSS.n11 0.0944005
R46 VSS.n11 VSS.n10 0.0944005
R47 VSS.n1 VSS.n0 0.0944005
R48 VSS.n4 VSS.n3 0.0944005
R49 VSS.n3 VSS.n2 0.0944005
R50 VSS.n7 VSS.n6 0.0640462
R51 VSS.n17 VSS.n16 0.0639407
R52 VSS.n21 VSS.n20 0.0591735
R53 VSS.t2 VSS.n7 0.0472599
R54 VSS.t0 VSS.n17 0.0471159
R55 VSS.n18 VSS.t0 0.0039133
R56 VSS.n8 VSS.t2 0.0039133
R57 VSS.n9 VSS.n8 0.0039133
R58 VSS.n19 VSS.n18 0.0039133
R59 VSS.n20 VSS.n19 0.00233287
R60 A.n0 A.t0 155.132
R61 A.n0 A.t1 140.864
R62 A A.n0 0.428385
C0 A VDD 0.266f
C1 OUT VDD 0.525f
C2 VDD B 0.266f
C3 OUT A 0.0821f
C4 A B 0.0265f
C5 VDD a_704_16# 0.00823f
C6 OUT B 0.297f
C7 A a_704_16# 0.0121f
C8 OUT a_704_16# 0.108f
C9 B a_704_16# 0.0121f
.ends

