* NGSPICE file created from inverter.ext - technology: sky130A

.subckt inverter Vin Vout VDD VSS
X0 Vout Vin.t1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1 Vout Vin.t0 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
R0 Vin.n0 Vin.t0 222.611
R1 Vin Vin.t1 140.625
R2 Vin.n0 Vin 0.6255
R3 Vin Vin.n0 0.038
R4 VDD.n7 VDD.n1 134.024
R5 VDD.n10 VDD.n7 106.049
R6 VDD.n12 VDD.n11 9.3005
R7 VDD VDD.n12 0.148
R8 VDD.n12 VDD.n10 0.117644
R9 VDD.n1 VDD.n0 0.0349892
R10 VDD.n3 VDD.n2 0.018623
R11 VDD.n7 VDD.n6 0.018623
R12 VDD.n4 VDD.n3 0.0140831
R13 VDD.n6 VDD.n5 0.0140829
R14 VDD.n5 VDD.n4 0.0115798
R15 VDD.n9 VDD.n8 0.00380159
R16 VDD.n10 VDD.n9 0.00142302
R17 VSS.n12 VSS.n9 116.329
R18 VSS.n5 VSS.n4 90.2269
R19 VSS.n13 VSS.n12 81.0463
R20 VSS.n14 VSS.n13 9.3005
R21 VSS VSS.n14 0.152286
R22 VSS.n14 VSS.n7 0.11402
R23 VSS.n9 VSS.n8 0.10956
R24 VSS.n12 VSS.n11 0.0944005
R25 VSS.n4 VSS.n3 0.0944005
R26 VSS.n11 VSS.n10 0.0485732
R27 VSS.n3 VSS.n2 0.0485718
R28 VSS.n7 VSS.n5 0.00690386
R29 VSS.n1 VSS.n0 0.0039133
R30 VSS.n5 VSS.n1 0.00366545
R31 VSS.n7 VSS.n6 0.000572701
C0 Vout Vin 0.166f
C1 VDD Vin 0.25f
C2 Vout VDD 0.326f
.ends

