** sch_path: /foss/designs/test/inv.sch
*.subckt inv VDD VSS IN OUT
*.ipin VDD
*.ipin VSS
*.ipin IN
*.opin OUT
XM1 OUT IN VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad=(int((nf+1)/2)*W/nf*0.29) as=(int((nf+2)/2)*W/nf*0.29)
+ pd=(2*int((nf+1)/2)*(W/nf+0.29)) ps=(2*int((nf+2)/2)*(W/nf+0.29)) nrd=(0.29/W) nrs=(0.29/W)
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 ad=(int((nf+1)/2)*W/nf*0.29) as=(int((nf+2)/2)*W/nf*0.29)
+ pd=(2*int((nf+1)/2)*(W/nf+0.29)) ps=(2*int((nf+2)/2)*(W/nf+0.29)) nrd=(0.29/W) nrs=(0.29/W)
+ sa=0 sb=0 sd=0 mult=1 m=1
*.ends
*.end
