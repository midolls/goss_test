magic
tech sky130A
magscale 1 2
timestamp 1691223565
<< error_p >>
rect -29 165 29 171
rect -29 131 -17 165
rect -29 125 29 131
rect -29 -131 29 -125
rect -29 -165 -17 -131
rect -29 -171 29 -165
<< nwell >>
rect -211 -303 211 303
<< pmos >>
rect -15 -84 15 84
<< pdiff >>
rect -73 72 -15 84
rect -73 -72 -61 72
rect -27 -72 -15 72
rect -73 -84 -15 -72
rect 15 72 73 84
rect 15 -72 27 72
rect 61 -72 73 72
rect 15 -84 73 -72
<< pdiffc >>
rect -61 -72 -27 72
rect 27 -72 61 72
<< nsubdiff >>
rect -175 233 -79 267
rect 79 233 175 267
rect -175 171 -141 233
rect 141 171 175 233
rect -175 -233 -141 -171
rect 141 -233 175 -171
rect -175 -267 -79 -233
rect 79 -267 175 -233
<< nsubdiffcont >>
rect -79 233 79 267
rect -175 -171 -141 171
rect 141 -171 175 171
rect -79 -267 79 -233
<< poly >>
rect -33 165 33 181
rect -33 131 -17 165
rect 17 131 33 165
rect -33 115 33 131
rect -15 84 15 115
rect -15 -115 15 -84
rect -33 -131 33 -115
rect -33 -165 -17 -131
rect 17 -165 33 -131
rect -33 -181 33 -165
<< polycont >>
rect -17 131 17 165
rect -17 -165 17 -131
<< locali >>
rect -175 233 -79 267
rect 79 233 175 267
rect -175 171 -141 233
rect 141 171 175 233
rect -33 131 -17 165
rect 17 131 33 165
rect -61 72 -27 88
rect -61 -88 -27 -72
rect 27 72 61 88
rect 27 -88 61 -72
rect -33 -165 -17 -131
rect 17 -165 33 -131
rect -175 -233 -141 -171
rect 141 -233 175 -171
rect -175 -267 -79 -233
rect 79 -267 175 -233
<< viali >>
rect -17 131 17 165
rect -61 -72 -27 72
rect 27 -72 61 72
rect -17 -165 17 -131
<< metal1 >>
rect -29 165 29 171
rect -29 131 -17 165
rect 17 131 29 165
rect -29 125 29 131
rect -67 72 -21 84
rect -67 -72 -61 72
rect -27 -72 -21 72
rect -67 -84 -21 -72
rect 21 72 67 84
rect 21 -72 27 72
rect 61 -72 67 72
rect 21 -84 67 -72
rect -29 -131 29 -125
rect -29 -165 -17 -131
rect 17 -165 29 -131
rect -29 -171 29 -165
<< properties >>
string FIXED_BBOX -158 -250 158 250
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.84 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
