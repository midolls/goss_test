* NGSPICE file created from ringosil.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_L78EGD a_n33_33# a_15_n73# a_n73_n73# a_n175_n185#
X0 a_15_n73# a_n33_33# a_n73_n73# a_n175_n185# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
C0 a_n73_n73# a_15_n73# 0.0699f
C1 a_15_n73# a_n33_33# 0.0121f
C2 a_n73_n73# a_n33_33# 0.0121f
C3 a_15_n73# a_n175_n185# 0.0789f
C4 a_n73_n73# a_n175_n185# 0.0789f
C5 a_n33_33# a_n175_n185# 0.221f
.ends

.subckt sky130_fd_pr__pfet_01v8_2ZD9BZ w_n211_n226# a_n73_n6# a_15_n6# a_n33_n103#
+ VSUBS
X0 a_15_n6# a_n33_n103# a_n73_n6# w_n211_n226# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
C0 w_n211_n226# a_15_n6# 0.0505f
C1 w_n211_n226# a_n33_n103# 0.146f
C2 a_n33_n103# a_15_n6# 0.0112f
C3 w_n211_n226# a_n73_n6# 0.0505f
C4 a_n73_n6# a_15_n6# 0.0699f
C5 a_n73_n6# a_n33_n103# 0.0112f
C6 a_15_n6# VSUBS 0.0283f
C7 a_n73_n6# VSUBS 0.0283f
C8 a_n33_n103# VSUBS 0.0809f
C9 w_n211_n226# VSUBS 0.899f
.ends

.subckt nand OUT VDD m1_1070_58# m1_670_62# m1_726_n34# VSS
Xsky130_fd_pr__nfet_01v8_L78EGD_0 m1_1070_58# OUT m1_726_n34# VSS sky130_fd_pr__nfet_01v8_L78EGD
XXM2 VDD VDD OUT m1_1070_58# VSS sky130_fd_pr__pfet_01v8_2ZD9BZ
XXM4 m1_670_62# m1_726_n34# VSS VSS sky130_fd_pr__nfet_01v8_L78EGD
Xsky130_fd_pr__pfet_01v8_2ZD9BZ_0 VDD VDD OUT m1_670_62# VSS sky130_fd_pr__pfet_01v8_2ZD9BZ
C0 VDD m1_670_62# 0.0497f
C1 m1_1070_58# m1_726_n34# 4.48e-19
C2 OUT m1_726_n34# 0.0302f
C3 m1_1070_58# OUT 0.225f
C4 m1_726_n34# m1_670_62# 1.78e-20
C5 m1_1070_58# m1_670_62# 0.0367f
C6 OUT m1_670_62# 0.0661f
C7 VDD m1_726_n34# 0.00668f
C8 VDD m1_1070_58# 0.0499f
C9 VDD OUT 0.31f
C10 m1_726_n34# VSS 0.307f
C11 m1_670_62# VSS 0.376f
C12 OUT VSS 0.455f
C13 m1_1070_58# VSS 0.318f
C14 VDD VSS 1.88f
.ends

.subckt sky130_fd_pr__pfet_01v8_2MG8BZ a_n73_n48# a_n33_n145# a_15_n48# w_n211_n268#
+ VSUBS
X0 a_15_n48# a_n33_n145# a_n73_n48# w_n211_n268# sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
C0 a_n33_n145# a_15_n48# 0.0137f
C1 w_n211_n268# a_15_n48# 0.0761f
C2 a_n73_n48# a_15_n48# 0.137f
C3 w_n211_n268# a_n33_n145# 0.144f
C4 a_n73_n48# a_n33_n145# 0.0137f
C5 a_n73_n48# w_n211_n268# 0.0761f
C6 a_15_n48# VSUBS 0.0453f
C7 a_n73_n48# VSUBS 0.0453f
C8 a_n33_n145# VSUBS 0.0804f
C9 w_n211_n268# VSUBS 1.05f
.ends

.subckt sky130_fd_pr__nfet_01v8_EDL9KC a_n33_33# a_15_n73# a_n73_n73# a_n175_n185#
X0 a_15_n73# a_n33_33# a_n73_n73# a_n175_n185# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
C0 a_n33_33# a_n73_n73# 0.0121f
C1 a_15_n73# a_n73_n73# 0.0699f
C2 a_15_n73# a_n33_33# 0.0121f
C3 a_15_n73# a_n175_n185# 0.0789f
C4 a_n73_n73# a_n175_n185# 0.0789f
C5 a_n33_33# a_n175_n185# 0.221f
.ends

.subckt inverter VDD Vin Vout VSS
Xsky130_fd_pr__pfet_01v8_2MG8BZ_0 VDD Vin Vout VDD VSS sky130_fd_pr__pfet_01v8_2MG8BZ
Xsky130_fd_pr__nfet_01v8_EDL9KC_0 Vin Vout VSS VSS sky130_fd_pr__nfet_01v8_EDL9KC
C0 Vin Vout 0.14f
C1 VDD Vout 0.113f
C2 VDD Vin 0.0921f
C3 Vout VSS 0.303f
C4 Vin VSS 0.382f
C5 VDD VSS 1.23f
.ends

.subckt ringosil VSS EN CLK VDD
Xx1 x2/Vin VDD CLK EN x1/m1_726_n34# VSS nand
Xx3 VDD x3/Vin x4/Vin VSS inverter
Xx2 VDD x2/Vin x3/Vin VSS inverter
Xx4 VDD x4/Vin x5/Vin VSS inverter
Xx5 VDD x5/Vin x6/Vin VSS inverter
Xx6 VDD x6/Vin x7/Vin VSS inverter
Xx7 VDD x7/Vin x8/Vin VSS inverter
Xx8 VDD x8/Vin x9/Vin VSS inverter
Xx9 VDD x9/Vin x9/Vout VSS inverter
Xx10 VDD x9/Vout x11/Vin VSS inverter
Xx11 VDD x11/Vin CLK VSS inverter
X0 x1/m1_726_n34# EN.t0 VSS VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X1 x2/Vin EN.t1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
R0 VDD.n16 VDD.n15 163.06
R1 VDD.n144 VDD.n143 161.287
R2 VDD.n96 VDD.n95 159.516
R3 VDD.n64 VDD.n63 159.516
R4 VDD.n128 VDD.n127 157.744
R5 VDD.n112 VDD.n111 155.97
R6 VDD.n48 VDD.n47 155.97
R7 VDD.n32 VDD.n31 155.97
R8 VDD.n183 VDD.n175 118.213
R9 VDD.n183 VDD.n182 118.213
R10 VDD.n171 VDD.n163 118.213
R11 VDD.n171 VDD.n165 118.213
R12 VDD.n93 VDD.n92 98.7195
R13 VDD.n109 VDD.n108 98.7195
R14 VDD.n125 VDD.n124 98.7195
R15 VDD.n141 VDD.n140 98.7195
R16 VDD.n158 VDD.n157 98.7195
R17 VDD.n67 VDD.n66 98.7195
R18 VDD.n51 VDD.n50 98.7195
R19 VDD.n35 VDD.n34 98.7195
R20 VDD.n19 VDD.n18 98.7195
R21 VDD.n2 VDD.n1 98.7195
R22 VDD.n82 VDD.n81 98.7195
R23 VDD.n99 VDD.n98 98.7195
R24 VDD.n115 VDD.n114 98.7195
R25 VDD.n131 VDD.n130 98.7195
R26 VDD.n147 VDD.n146 98.7195
R27 VDD.n78 VDD.n77 98.7195
R28 VDD.n61 VDD.n60 98.7195
R29 VDD.n45 VDD.n44 98.7195
R30 VDD.n29 VDD.n28 98.7195
R31 VDD.n13 VDD.n12 98.7195
R32 VDD.n12 VDD.n11 9.3005
R33 VDD.n3 VDD.n2 9.3005
R34 VDD.n28 VDD.n27 9.3005
R35 VDD.n20 VDD.n19 9.3005
R36 VDD.n44 VDD.n43 9.3005
R37 VDD.n36 VDD.n35 9.3005
R38 VDD.n60 VDD.n59 9.3005
R39 VDD.n52 VDD.n51 9.3005
R40 VDD.n79 VDD.n78 9.3005
R41 VDD.n68 VDD.n67 9.3005
R42 VDD.n148 VDD.n147 9.3005
R43 VDD.n159 VDD.n158 9.3005
R44 VDD.n132 VDD.n131 9.3005
R45 VDD.n140 VDD.n139 9.3005
R46 VDD.n116 VDD.n115 9.3005
R47 VDD.n124 VDD.n123 9.3005
R48 VDD.n100 VDD.n99 9.3005
R49 VDD.n108 VDD.n107 9.3005
R50 VDD.n83 VDD.n82 9.3005
R51 VDD.n92 VDD.n91 9.3005
R52 VDD.n83 VDD.n79 3.56641
R53 VDD.n184 VDD.n172 0.515806
R54 VDD.n172 VDD 0.264531
R55 VDD VDD.n184 0.256878
R56 VDD.n68 VDD 0.148
R57 VDD.n52 VDD 0.148
R58 VDD.n36 VDD 0.148
R59 VDD.n20 VDD 0.148
R60 VDD.n3 VDD 0.148
R61 VDD.n91 VDD 0.148
R62 VDD.n107 VDD 0.148
R63 VDD.n123 VDD 0.148
R64 VDD.n139 VDD 0.148
R65 VDD.n160 VDD.n159 0.1355
R66 VDD.n11 VDD 0.1305
R67 VDD.n148 VDD 0.12925
R68 VDD.n59 VDD 0.128
R69 VDD.n100 VDD 0.128
R70 VDD.n132 VDD 0.12675
R71 VDD.n43 VDD 0.1255
R72 VDD.n27 VDD 0.1255
R73 VDD.n116 VDD 0.1255
R74 VDD.n79 VDD.n75 0.11675
R75 VDD.n75 VDD.n68 0.11675
R76 VDD.n59 VDD.n58 0.11675
R77 VDD.n58 VDD.n52 0.11675
R78 VDD.n43 VDD.n42 0.11675
R79 VDD.n42 VDD.n36 0.11675
R80 VDD.n27 VDD.n26 0.11675
R81 VDD.n26 VDD.n20 0.11675
R82 VDD.n11 VDD.n10 0.11675
R83 VDD.n10 VDD.n3 0.11675
R84 VDD.n90 VDD.n83 0.11675
R85 VDD.n91 VDD.n90 0.11675
R86 VDD.n106 VDD.n100 0.11675
R87 VDD.n107 VDD.n106 0.11675
R88 VDD.n122 VDD.n116 0.11675
R89 VDD.n123 VDD.n122 0.11675
R90 VDD.n138 VDD.n132 0.11675
R91 VDD.n139 VDD.n138 0.11675
R92 VDD.n154 VDD.n148 0.11675
R93 VDD.n159 VDD.n154 0.11675
R94 VDD.n167 VDD.n166 0.0349892
R95 VDD.n177 VDD.n176 0.0349892
R96 VDD.n178 VDD.n177 0.0349892
R97 VDD.n134 VDD.n133 0.0349892
R98 VDD.n135 VDD.n134 0.0349892
R99 VDD.n118 VDD.n117 0.0349892
R100 VDD.n119 VDD.n118 0.0349892
R101 VDD.n102 VDD.n101 0.0349892
R102 VDD.n103 VDD.n102 0.0349892
R103 VDD.n85 VDD.n84 0.0349892
R104 VDD.n150 VDD.n149 0.0349892
R105 VDD.n151 VDD.n150 0.0349892
R106 VDD.n22 VDD.n21 0.0349892
R107 VDD.n23 VDD.n22 0.0349892
R108 VDD.n38 VDD.n37 0.0349892
R109 VDD.n39 VDD.n38 0.0349892
R110 VDD.n54 VDD.n53 0.0349892
R111 VDD.n55 VDD.n54 0.0349892
R112 VDD.n70 VDD.n69 0.0349892
R113 VDD.n71 VDD.n70 0.0349892
R114 VDD.n5 VDD.n4 0.0349892
R115 VDD.n6 VDD.n5 0.0292476
R116 VDD.n86 VDD.n85 0.0292024
R117 VDD.n165 VDD.n164 0.0286326
R118 VDD.n163 VDD.n162 0.0286326
R119 VDD.n162 VDD.n161 0.0286326
R120 VDD.n182 VDD.n181 0.0286326
R121 VDD.n181 VDD.n180 0.0286326
R122 VDD.n175 VDD.n174 0.0286326
R123 VDD.n174 VDD.n173 0.0286326
R124 VDD.n168 VDD.n167 0.0275362
R125 VDD.n130 VDD.n129 0.018623
R126 VDD.n129 VDD.n128 0.018623
R127 VDD.n142 VDD.n141 0.018623
R128 VDD.n143 VDD.n142 0.018623
R129 VDD.n114 VDD.n113 0.018623
R130 VDD.n113 VDD.n112 0.018623
R131 VDD.n126 VDD.n125 0.018623
R132 VDD.n127 VDD.n126 0.018623
R133 VDD.n98 VDD.n97 0.018623
R134 VDD.n97 VDD.n96 0.018623
R135 VDD.n110 VDD.n109 0.018623
R136 VDD.n111 VDD.n110 0.018623
R137 VDD.n81 VDD.n80 0.018623
R138 VDD.n94 VDD.n93 0.018623
R139 VDD.n95 VDD.n94 0.018623
R140 VDD.n157 VDD.n156 0.018623
R141 VDD.n156 VDD.n155 0.018623
R142 VDD.n146 VDD.n145 0.018623
R143 VDD.n145 VDD.n144 0.018623
R144 VDD.n18 VDD.n17 0.018623
R145 VDD.n17 VDD.n16 0.018623
R146 VDD.n30 VDD.n29 0.018623
R147 VDD.n31 VDD.n30 0.018623
R148 VDD.n34 VDD.n33 0.018623
R149 VDD.n33 VDD.n32 0.018623
R150 VDD.n46 VDD.n45 0.018623
R151 VDD.n47 VDD.n46 0.018623
R152 VDD.n50 VDD.n49 0.018623
R153 VDD.n49 VDD.n48 0.018623
R154 VDD.n62 VDD.n61 0.018623
R155 VDD.n63 VDD.n62 0.018623
R156 VDD.n66 VDD.n65 0.018623
R157 VDD.n65 VDD.n64 0.018623
R158 VDD.n77 VDD.n76 0.018623
R159 VDD.n1 VDD.n0 0.018623
R160 VDD.n14 VDD.n13 0.018623
R161 VDD.n15 VDD.n14 0.018623
R162 VDD VDD.n160 0.0130883
R163 VDD.n160 VDD 0.013
R164 VDD.n169 VDD.n168 0.00895217
R165 VDD.n7 VDD.n6 0.00748901
R166 VDD.n87 VDD.n86 0.00728604
R167 VDD VDD 0.00560204
R168 VDD.n137 VDD.n136 0.00380159
R169 VDD.n136 VDD.n135 0.00380159
R170 VDD.n121 VDD.n120 0.00380159
R171 VDD.n120 VDD.n119 0.00380159
R172 VDD.n105 VDD.n104 0.00380159
R173 VDD.n104 VDD.n103 0.00380159
R174 VDD.n89 VDD.n88 0.00380159
R175 VDD.n88 VDD.n87 0.00380159
R176 VDD.n9 VDD.n8 0.00380159
R177 VDD.n8 VDD.n7 0.00380159
R178 VDD.n25 VDD.n24 0.00380159
R179 VDD.n24 VDD.n23 0.00380159
R180 VDD.n41 VDD.n40 0.00380159
R181 VDD.n40 VDD.n39 0.00380159
R182 VDD.n57 VDD.n56 0.00380159
R183 VDD.n56 VDD.n55 0.00380159
R184 VDD.n74 VDD.n73 0.00380159
R185 VDD.n153 VDD.n152 0.00380159
R186 VDD.n152 VDD.n151 0.00380159
R187 VDD.n183 VDD.n179 0.00380159
R188 VDD.n179 VDD.n178 0.00380159
R189 VDD.n171 VDD.n170 0.00380159
R190 VDD.n170 VDD.n169 0.00380159
R191 VDD.n73 VDD.n72 0.00369982
R192 VDD.n184 VDD.n183 0.00233287
R193 VDD.n172 VDD.n171 0.00233287
R194 VDD.n72 VDD.n71 0.00160176
R195 VDD.n10 VDD.n9 0.000567328
R196 VDD.n26 VDD.n25 0.000567328
R197 VDD.n42 VDD.n41 0.000567328
R198 VDD.n58 VDD.n57 0.000567328
R199 VDD.n75 VDD.n74 0.000567328
R200 VDD.n154 VDD.n153 0.000567328
R201 VDD.n138 VDD.n137 0.000567328
R202 VDD.n122 VDD.n121 0.000567328
R203 VDD.n106 VDD.n105 0.000567328
R204 VDD.n90 VDD.n89 0.000567328
R205 EN.n0 EN.t1 155.304
R206 EN.n0 EN.t0 140.912
R207 EN EN.n0 0.178234
C0 VDD x2/Vin 0.0529f
C1 x9/Vout x4/Vin 9.79e-20
C2 VDD x4/Vin 0.0569f
C3 x8/Vin x5/Vin 0.0031f
C4 VDD x6/Vin 0.0536f
C5 VDD x5/Vin 0.0568f
C6 x9/Vout x11/Vin 0.0163f
C7 VDD x11/Vin 0.052f
C8 x8/Vin x9/Vin 0.0179f
C9 VDD x1/m1_726_n34# -6.53e-20
C10 CLK EN 0.00189f
C11 x3/Vin x9/Vout 0.0031f
C12 x3/Vin VDD 0.0578f
C13 x9/Vout x9/Vin 0.018f
C14 VDD x9/Vin 0.0568f
C15 EN x2/Vin 0.00141f
C16 VDD x8/Vin 0.0605f
C17 x7/Vin x6/Vin 0.0111f
C18 VDD x9/Vout 0.0539f
C19 CLK x2/Vin 0.0643f
C20 CLK x4/Vin 6.89e-19
C21 x4/Vin x2/Vin 1.29e-19
C22 CLK x5/Vin 2.81e-19
C23 x6/Vin x2/Vin 1.23e-20
C24 CLK x11/Vin 0.0106f
C25 x5/Vin x2/Vin 5.75e-20
C26 x4/Vin x5/Vin 0.018f
C27 x2/Vin x11/Vin 0.0031f
C28 x6/Vin x5/Vin 0.0179f
C29 VDD EN 0.0142f
C30 CLK x1/m1_726_n34# 0.0278f
C31 x3/Vin CLK 0.00525f
C32 x7/Vin x8/Vin 0.014f
C33 CLK x9/Vin 5e-19
C34 x1/m1_726_n34# x2/Vin -9.89e-20
C35 x3/Vin x2/Vin 0.0126f
C36 x7/Vin VDD 0.601f
C37 x3/Vin x4/Vin 0.0179f
C38 x4/Vin x9/Vin 0.0031f
C39 x8/Vin CLK 8.14e-20
C40 x3/Vin x11/Vin 9.79e-20
C41 x9/Vin x5/Vin 9.41e-20
C42 x9/Vout CLK 0.00103f
C43 VDD CLK 0.0322f
C44 x8/Vin x6/Vin 9.41e-20
C45 x11/Vin VSS 0.35f
C46 x9/Vout VSS 0.34f
C47 x9/Vin VSS 0.334f
C48 x8/Vin VSS 0.335f
C49 x7/Vin VSS 0.605f
C50 x6/Vin VSS 0.349f
C51 x5/Vin VSS 0.334f
C52 x4/Vin VSS 0.334f
C53 x3/Vin VSS 0.338f
C54 x1/m1_726_n34# VSS 0.137f
C55 EN VSS 0.357f
C56 x2/Vin VSS 0.545f
C57 CLK VSS 0.953f
C58 VDD VSS 11.2f
.ends

