* NGSPICE file created from inv.ext - technology: sky130A

.subckt inv IN OUT VDD VSS
X0 OUT.t0 IN.t0 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X1 OUT.t1 IN.t1 VSS.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
R0 IN.n0 IN.t0 222.768
R1 IN.n0 IN.t1 140.803
R2 IN IN.n0 0.827706
R3 VDD.n9 VDD.n8 134.024
R4 VDD.n9 VDD.n1 134.024
R5 VDD.n10 VDD.t1 34.4686
R6 VDD VDD.n11 1.05428
R7 VDD.n10 VDD 0.243233
R8 VDD.n11 VDD.n10 0.0644535
R9 VDD.n3 VDD.n2 0.0349892
R10 VDD.t0 VDD.n3 0.0349892
R11 VDD.n8 VDD.n7 0.018623
R12 VDD.n1 VDD.n0 0.018623
R13 VDD.t0 VDD.n4 0.0135718
R14 VDD.n6 VDD.n5 0.00383554
R15 VDD.n9 VDD.n6 0.00380159
R16 VDD.n11 VDD.n9 0.00233287
R17 VDD.n5 VDD.t0 0.00163201
R18 OUT OUT.t1 42.4221
R19 OUT OUT.t0 35.1823
R20 VSS.n9 VSS.n1 116.329
R21 VSS.n9 VSS.n8 116.329
R22 VSS.n10 VSS.t1 41.7438
R23 VSS VSS.n10 0.244686
R24 VSS.n3 VSS.n2 0.10956
R25 VSS.n1 VSS.n0 0.0944005
R26 VSS.n8 VSS.n7 0.0944005
R27 VSS.n10 VSS.n9 0.0648329
R28 VSS.n4 VSS.n3 0.0591703
R29 VSS.t0 VSS.n4 0.052136
R30 VSS.n9 VSS.n6 0.0039133
R31 VSS.n6 VSS.n5 0.00281698
R32 VSS.n5 VSS.t0 0.00259631
C0 VDD IN 0.248f
C1 OUT VDD 0.322f
C2 OUT IN 0.144f
.ends

