* NGSPICE file created from ringosil.ext - technology: sky130A

.subckt ringosil EN CLK VDD VSS
X0 x7.Vin x6.Vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X1 VDD x11.Vin CLK VDD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X2 x2/Vin CLK.t1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X3 x5.Vin x4.Vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X4 x6.Vin x5.Vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X5 VDD x9.Vout x11.Vin VDD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X6 x3.Vin x2.Vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X7 VDD x9.Vin x9.Vout VDD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X8 VDD x7.Vin x8.Vin VDD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X9 x4.Vin x3.Vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X10 x2/Vin EN.t1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X11 x2/Vin CLK.t0 x1/m1_726_n34# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X12 VDD x8.Vin x9.Vin VDD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
R0 CLK.n0 CLK.t1 155.758
R1 CLK.n0 CLK.t0 140.583
R2 CLK CLK.n0 4.52884
R3 x11/Vout CLK 0.438
R4 VSS.n19 VSS.n16 64770.9
R5 VSS.n16 VSS.n15 49622.2
R6 VSS.n14 VSS.n13 49500
R7 VSS.n15 VSS.n14 49377.8
R8 VSS.n45 VSS.n44 263.205
R9 VSS.n75 VSS.n74 263.205
R10 VSS.n105 VSS.n104 263.205
R11 VSS.n138 VSS.n137 263.205
R12 VSS.n191 VSS.n190 218.511
R13 VSS.n141 VSS.n138 188.714
R14 VSS.n48 VSS.n45 183.748
R15 VSS.n78 VSS.n75 173.815
R16 VSS.n106 VSS.n105 173.815
R17 VSS.n194 VSS.n185 116.329
R18 VSS.n194 VSS.n193 116.329
R19 VSS.n181 VSS.n173 116.329
R20 VSS.n181 VSS.n180 116.329
R21 VSS.n114 VSS.n113 82.9914
R22 VSS.n11 VSS.n10 82.6358
R23 VSS.n8 VSS.n7 82.6358
R24 VSS.n5 VSS.n4 82.6358
R25 VSS.n1 VSS.n0 82.6358
R26 VSS.n22 VSS.n21 81.4018
R27 VSS.n51 VSS.n50 81.4018
R28 VSS.n81 VSS.n80 81.4018
R29 VSS.n109 VSS.n108 81.4018
R30 VSS.n144 VSS.n143 81.4018
R31 VSS.n135 VSS.n134 81.0463
R32 VSS.n102 VSS.n101 81.0463
R33 VSS.n72 VSS.n71 81.0463
R34 VSS.n42 VSS.n41 81.0463
R35 VSS.n169 VSS.n168 81.0463
R36 VSS.n24 VSS.n22 9.30308
R37 VSS.n170 VSS.n169 9.3005
R38 VSS.n147 VSS.n146 9.3005
R39 VSS.n145 VSS.n144 9.3005
R40 VSS.n163 VSS.n162 9.3005
R41 VSS.n110 VSS.n109 9.3005
R42 VSS.n82 VSS.n81 9.3005
R43 VSS.n52 VSS.n51 9.3005
R44 VSS.n24 VSS.n23 9.3005
R45 VSS.n41 VSS.n40 9.3005
R46 VSS.n54 VSS.n53 9.3005
R47 VSS.n71 VSS.n70 9.3005
R48 VSS.n84 VSS.n83 9.3005
R49 VSS.n101 VSS.n100 9.3005
R50 VSS.n115 VSS.n114 9.3005
R51 VSS.n134 VSS.n133 9.3005
R52 VSS.n137 VSS.n3 4.96664
R53 x11/VSS x1/VSS 0.522407
R54 VSS.n195 VSS.n182 0.515806
R55 VSS.n182 x1/VSS 0.254327
R56 x11/VSS VSS.n195 0.249224
R57 VSS.n175 VSS.n174 0.10956
R58 VSS.n187 VSS.n186 0.10956
R59 VSS.n188 VSS.n187 0.10956
R60 VSS.n155 VSS.n154 0.10956
R61 VSS.n156 VSS.n155 0.10956
R62 VSS.n119 VSS.n118 0.10956
R63 VSS.n120 VSS.n119 0.10956
R64 VSS.n88 VSS.n87 0.10956
R65 VSS.n91 VSS.n88 0.10956
R66 VSS.n58 VSS.n57 0.10956
R67 VSS.n61 VSS.n58 0.10956
R68 VSS.n28 VSS.n27 0.10956
R69 VSS.n31 VSS.n28 0.10956
R70 VSS.n30 VSS.n29 0.10956
R71 VSS.n31 VSS.n30 0.10956
R72 VSS.n60 VSS.n59 0.10956
R73 VSS.n61 VSS.n60 0.10956
R74 VSS.n90 VSS.n89 0.10956
R75 VSS.n91 VSS.n90 0.10956
R76 VSS.n125 VSS.n124 0.10956
R77 VSS.n126 VSS.n125 0.10956
R78 VSS.n153 VSS.n152 0.10956
R79 VSS.n156 VSS.n153 0.10956
R80 VSS.n180 VSS.n179 0.0944005
R81 VSS.n173 VSS.n172 0.0944005
R82 VSS.n172 VSS.n171 0.0944005
R83 VSS.n193 VSS.n192 0.0944005
R84 VSS.n192 VSS.n191 0.0944005
R85 VSS.n185 VSS.n184 0.0944005
R86 VSS.n184 VSS.n183 0.0944005
R87 VSS.n143 VSS.n142 0.0944005
R88 VSS.n142 VSS.n141 0.0944005
R89 VSS.n165 VSS.n164 0.0944005
R90 VSS.n166 VSS.n165 0.0944005
R91 VSS.n108 VSS.n107 0.0944005
R92 VSS.n107 VSS.n106 0.0944005
R93 VSS.n2 VSS.n1 0.0944005
R94 VSS.n3 VSS.n2 0.0944005
R95 VSS.n80 VSS.n79 0.0944005
R96 VSS.n79 VSS.n78 0.0944005
R97 VSS.n6 VSS.n5 0.0944005
R98 VSS.n104 VSS.n6 0.0944005
R99 VSS.n50 VSS.n49 0.0944005
R100 VSS.n49 VSS.n48 0.0944005
R101 VSS.n9 VSS.n8 0.0944005
R102 VSS.n74 VSS.n9 0.0944005
R103 VSS.n21 VSS.n20 0.0944005
R104 VSS.n20 VSS.n19 0.0944005
R105 VSS.n12 VSS.n11 0.0944005
R106 VSS.n44 VSS.n12 0.0944005
R107 VSS.n18 VSS.n17 0.0944005
R108 VSS.n19 VSS.n18 0.0944005
R109 VSS.n43 VSS.n42 0.0944005
R110 VSS.n44 VSS.n43 0.0944005
R111 VSS.n47 VSS.n46 0.0944005
R112 VSS.n48 VSS.n47 0.0944005
R113 VSS.n73 VSS.n72 0.0944005
R114 VSS.n74 VSS.n73 0.0944005
R115 VSS.n77 VSS.n76 0.0944005
R116 VSS.n78 VSS.n77 0.0944005
R117 VSS.n103 VSS.n102 0.0944005
R118 VSS.n104 VSS.n103 0.0944005
R119 VSS.n113 VSS.n112 0.0944005
R120 VSS.n112 VSS.n111 0.0944005
R121 VSS.n136 VSS.n135 0.0944005
R122 VSS.n137 VSS.n136 0.0944005
R123 VSS.n168 VSS.n167 0.0944005
R124 VSS.n167 VSS.n166 0.0944005
R125 VSS.n140 VSS.n139 0.0944005
R126 VSS.n141 VSS.n140 0.0944005
R127 VSS.n40 x7/VSS 0.0771753
R128 VSS.n70 x5/VSS 0.0771753
R129 VSS.n100 x9/VSS 0.0771753
R130 x11/VSS VSS.n170 0.0771753
R131 VSS.n176 VSS.n175 0.0768221
R132 VSS.n133 x10/VSS 0.0765309
R133 VSS.n145 x3/VSS 0.066866
R134 VSS.n52 x7/VSS 0.0662216
R135 VSS.n82 x5/VSS 0.064933
R136 VSS.n110 x9/VSS 0.064933
R137 VSS.n39 VSS.n38 0.055268
R138 VSS.n69 VSS.n68 0.055268
R139 VSS.n99 VSS.n98 0.055268
R140 VSS.n163 VSS.n161 0.055268
R141 VSS.n26 VSS.n24 0.0546237
R142 VSS.n56 VSS.n54 0.0546237
R143 VSS.n86 VSS.n84 0.0546237
R144 VSS.n132 VSS.n131 0.0546237
R145 VSS.n149 VSS.n147 0.0546237
R146 VSS.n117 VSS.n115 0.0539794
R147 VSS.n177 VSS.n176 0.0342337
R148 VSS.n159 VSS.n151 0.00396756
R149 VSS.n123 VSS.n122 0.00396756
R150 VSS.n96 VSS.n93 0.00396756
R151 VSS.n66 VSS.n63 0.00396756
R152 VSS.n36 VSS.n33 0.00396756
R153 VSS.n36 VSS.n35 0.00396756
R154 VSS.n66 VSS.n65 0.00396756
R155 VSS.n96 VSS.n95 0.00396756
R156 VSS.n129 VSS.n128 0.00396756
R157 VSS.n159 VSS.n158 0.00396756
R158 VSS.n151 VSS.n150 0.0039133
R159 VSS.n122 VSS.n121 0.0039133
R160 VSS.n121 VSS.n120 0.0039133
R161 VSS.n93 VSS.n92 0.0039133
R162 VSS.n92 VSS.n91 0.0039133
R163 VSS.n63 VSS.n62 0.0039133
R164 VSS.n62 VSS.n61 0.0039133
R165 VSS.n33 VSS.n32 0.0039133
R166 VSS.n32 VSS.n31 0.0039133
R167 VSS.n35 VSS.n34 0.0039133
R168 VSS.n65 VSS.n64 0.0039133
R169 VSS.n95 VSS.n94 0.0039133
R170 VSS.n128 VSS.n127 0.0039133
R171 VSS.n127 VSS.n126 0.0039133
R172 VSS.n158 VSS.n157 0.0039133
R173 VSS.n157 VSS.n156 0.0039133
R174 VSS.n181 VSS.n178 0.0039133
R175 VSS.n178 VSS.n177 0.0039133
R176 VSS.n194 VSS.n189 0.0039133
R177 VSS.n189 VSS.n188 0.0039133
R178 VSS.n115 VSS.n110 0.00372165
R179 VSS.n133 VSS.n132 0.00372165
R180 VSS.n36 VSS.n26 0.00307732
R181 VSS.n38 VSS.n36 0.00307732
R182 VSS.n40 VSS.n39 0.00307732
R183 VSS.n54 VSS.n52 0.00307732
R184 VSS.n66 VSS.n56 0.00307732
R185 VSS.n68 VSS.n66 0.00307732
R186 VSS.n70 VSS.n69 0.00307732
R187 VSS.n84 VSS.n82 0.00307732
R188 VSS.n96 VSS.n86 0.00307732
R189 VSS.n98 VSS.n96 0.00307732
R190 VSS.n100 VSS.n99 0.00307732
R191 VSS.n123 VSS.n117 0.00307732
R192 VSS.n131 VSS.n129 0.00307732
R193 VSS.n147 VSS.n145 0.00307732
R194 VSS.n159 VSS.n149 0.00307732
R195 VSS.n161 VSS.n159 0.00307732
R196 VSS.n170 VSS.n163 0.00307732
R197 VSS.n182 VSS.n181 0.00233287
R198 VSS.n195 VSS.n194 0.00233287
R199 VSS.n129 VSS.n123 0.00114433
R200 x10/VSS x3/VSS 0.00114433
R201 VSS.n161 VSS.n160 0.000572701
R202 VSS.n149 VSS.n148 0.000572701
R203 VSS.n117 VSS.n116 0.000572701
R204 VSS.n86 VSS.n85 0.000572701
R205 VSS.n56 VSS.n55 0.000572701
R206 VSS.n26 VSS.n25 0.000572701
R207 VSS.n38 VSS.n37 0.000572701
R208 VSS.n68 VSS.n67 0.000572701
R209 VSS.n98 VSS.n97 0.000572701
R210 VSS.n131 VSS.n130 0.000572701
R211 VDD.n16 VDD.n15 163.06
R212 VDD.n144 VDD.n143 161.287
R213 VDD.n96 VDD.n95 159.516
R214 VDD.n64 VDD.n63 159.516
R215 VDD.n128 VDD.n127 157.744
R216 VDD.n112 VDD.n111 155.97
R217 VDD.n48 VDD.n47 155.97
R218 VDD.n32 VDD.n31 155.97
R219 VDD.n183 VDD.n175 118.213
R220 VDD.n183 VDD.n182 118.213
R221 VDD.n171 VDD.n163 118.213
R222 VDD.n171 VDD.n165 118.213
R223 VDD.n93 VDD.n92 98.7195
R224 VDD.n109 VDD.n108 98.7195
R225 VDD.n125 VDD.n124 98.7195
R226 VDD.n141 VDD.n140 98.7195
R227 VDD.n158 VDD.n157 98.7195
R228 VDD.n67 VDD.n66 98.7195
R229 VDD.n51 VDD.n50 98.7195
R230 VDD.n35 VDD.n34 98.7195
R231 VDD.n19 VDD.n18 98.7195
R232 VDD.n2 VDD.n1 98.7195
R233 VDD.n82 VDD.n81 98.7195
R234 VDD.n99 VDD.n98 98.7195
R235 VDD.n115 VDD.n114 98.7195
R236 VDD.n131 VDD.n130 98.7195
R237 VDD.n147 VDD.n146 98.7195
R238 VDD.n78 VDD.n77 98.7195
R239 VDD.n61 VDD.n60 98.7195
R240 VDD.n45 VDD.n44 98.7195
R241 VDD.n29 VDD.n28 98.7195
R242 VDD.n13 VDD.n12 98.7195
R243 VDD.n12 VDD.n11 9.3005
R244 VDD.n3 VDD.n2 9.3005
R245 VDD.n28 VDD.n27 9.3005
R246 VDD.n20 VDD.n19 9.3005
R247 VDD.n44 VDD.n43 9.3005
R248 VDD.n36 VDD.n35 9.3005
R249 VDD.n60 VDD.n59 9.3005
R250 VDD.n52 VDD.n51 9.3005
R251 VDD.n79 VDD.n78 9.3005
R252 VDD.n68 VDD.n67 9.3005
R253 VDD.n148 VDD.n147 9.3005
R254 VDD.n159 VDD.n158 9.3005
R255 VDD.n132 VDD.n131 9.3005
R256 VDD.n140 VDD.n139 9.3005
R257 VDD.n116 VDD.n115 9.3005
R258 VDD.n124 VDD.n123 9.3005
R259 VDD.n100 VDD.n99 9.3005
R260 VDD.n108 VDD.n107 9.3005
R261 VDD.n83 VDD.n82 9.3005
R262 VDD.n92 VDD.n91 9.3005
R263 VDD.n83 VDD.n79 3.56641
R264 VDD.n184 VDD.n172 0.515806
R265 VDD.n172 VDD 0.264531
R266 x2/VDD VDD.n184 0.256878
R267 VDD.n68 x7/VDD 0.148
R268 VDD.n52 x8/VDD 0.148
R269 VDD.n36 x9/VDD 0.148
R270 VDD.n20 x10/VDD 0.148
R271 VDD.n3 x11/VDD 0.148
R272 VDD.n91 x6/VDD 0.148
R273 VDD.n107 x5/VDD 0.148
R274 VDD.n123 x4/VDD 0.148
R275 VDD.n139 x3/VDD 0.148
R276 VDD.n160 VDD.n159 0.1355
R277 VDD.n11 x10/VDD 0.1305
R278 VDD.n148 x3/VDD 0.12925
R279 VDD.n59 x7/VDD 0.128
R280 VDD.n100 x6/VDD 0.128
R281 VDD.n132 x4/VDD 0.12675
R282 VDD.n43 x8/VDD 0.1255
R283 VDD.n27 x9/VDD 0.1255
R284 VDD.n116 x5/VDD 0.1255
R285 VDD.n79 VDD.n75 0.11675
R286 VDD.n75 VDD.n68 0.11675
R287 VDD.n59 VDD.n58 0.11675
R288 VDD.n58 VDD.n52 0.11675
R289 VDD.n43 VDD.n42 0.11675
R290 VDD.n42 VDD.n36 0.11675
R291 VDD.n27 VDD.n26 0.11675
R292 VDD.n26 VDD.n20 0.11675
R293 VDD.n11 VDD.n10 0.11675
R294 VDD.n10 VDD.n3 0.11675
R295 VDD.n90 VDD.n83 0.11675
R296 VDD.n91 VDD.n90 0.11675
R297 VDD.n106 VDD.n100 0.11675
R298 VDD.n107 VDD.n106 0.11675
R299 VDD.n122 VDD.n116 0.11675
R300 VDD.n123 VDD.n122 0.11675
R301 VDD.n138 VDD.n132 0.11675
R302 VDD.n139 VDD.n138 0.11675
R303 VDD.n154 VDD.n148 0.11675
R304 VDD.n159 VDD.n154 0.11675
R305 VDD.n167 VDD.n166 0.0349892
R306 VDD.n177 VDD.n176 0.0349892
R307 VDD.n178 VDD.n177 0.0349892
R308 VDD.n134 VDD.n133 0.0349892
R309 VDD.n135 VDD.n134 0.0349892
R310 VDD.n118 VDD.n117 0.0349892
R311 VDD.n119 VDD.n118 0.0349892
R312 VDD.n102 VDD.n101 0.0349892
R313 VDD.n103 VDD.n102 0.0349892
R314 VDD.n85 VDD.n84 0.0349892
R315 VDD.n150 VDD.n149 0.0349892
R316 VDD.n151 VDD.n150 0.0349892
R317 VDD.n22 VDD.n21 0.0349892
R318 VDD.n23 VDD.n22 0.0349892
R319 VDD.n38 VDD.n37 0.0349892
R320 VDD.n39 VDD.n38 0.0349892
R321 VDD.n54 VDD.n53 0.0349892
R322 VDD.n55 VDD.n54 0.0349892
R323 VDD.n70 VDD.n69 0.0349892
R324 VDD.n71 VDD.n70 0.0349892
R325 VDD.n5 VDD.n4 0.0349892
R326 VDD.n6 VDD.n5 0.0292476
R327 VDD.n86 VDD.n85 0.0292024
R328 VDD.n165 VDD.n164 0.0286326
R329 VDD.n163 VDD.n162 0.0286326
R330 VDD.n162 VDD.n161 0.0286326
R331 VDD.n182 VDD.n181 0.0286326
R332 VDD.n181 VDD.n180 0.0286326
R333 VDD.n175 VDD.n174 0.0286326
R334 VDD.n174 VDD.n173 0.0286326
R335 VDD.n168 VDD.n167 0.0275362
R336 VDD.n130 VDD.n129 0.018623
R337 VDD.n129 VDD.n128 0.018623
R338 VDD.n142 VDD.n141 0.018623
R339 VDD.n143 VDD.n142 0.018623
R340 VDD.n114 VDD.n113 0.018623
R341 VDD.n113 VDD.n112 0.018623
R342 VDD.n126 VDD.n125 0.018623
R343 VDD.n127 VDD.n126 0.018623
R344 VDD.n98 VDD.n97 0.018623
R345 VDD.n97 VDD.n96 0.018623
R346 VDD.n110 VDD.n109 0.018623
R347 VDD.n111 VDD.n110 0.018623
R348 VDD.n81 VDD.n80 0.018623
R349 VDD.n94 VDD.n93 0.018623
R350 VDD.n95 VDD.n94 0.018623
R351 VDD.n157 VDD.n156 0.018623
R352 VDD.n156 VDD.n155 0.018623
R353 VDD.n146 VDD.n145 0.018623
R354 VDD.n145 VDD.n144 0.018623
R355 VDD.n18 VDD.n17 0.018623
R356 VDD.n17 VDD.n16 0.018623
R357 VDD.n30 VDD.n29 0.018623
R358 VDD.n31 VDD.n30 0.018623
R359 VDD.n34 VDD.n33 0.018623
R360 VDD.n33 VDD.n32 0.018623
R361 VDD.n46 VDD.n45 0.018623
R362 VDD.n47 VDD.n46 0.018623
R363 VDD.n50 VDD.n49 0.018623
R364 VDD.n49 VDD.n48 0.018623
R365 VDD.n62 VDD.n61 0.018623
R366 VDD.n63 VDD.n62 0.018623
R367 VDD.n66 VDD.n65 0.018623
R368 VDD.n65 VDD.n64 0.018623
R369 VDD.n77 VDD.n76 0.018623
R370 VDD.n1 VDD.n0 0.018623
R371 VDD.n14 VDD.n13 0.018623
R372 VDD.n15 VDD.n14 0.018623
R373 x2/VDD VDD.n160 0.0130883
R374 VDD.n160 x2/VDD 0.013
R375 VDD.n169 VDD.n168 0.00895217
R376 VDD.n7 VDD.n6 0.00748901
R377 VDD.n87 VDD.n86 0.00728604
R378 VDD x1/VDD 0.00560204
R379 VDD.n137 VDD.n136 0.00380159
R380 VDD.n136 VDD.n135 0.00380159
R381 VDD.n121 VDD.n120 0.00380159
R382 VDD.n120 VDD.n119 0.00380159
R383 VDD.n105 VDD.n104 0.00380159
R384 VDD.n104 VDD.n103 0.00380159
R385 VDD.n89 VDD.n88 0.00380159
R386 VDD.n88 VDD.n87 0.00380159
R387 VDD.n9 VDD.n8 0.00380159
R388 VDD.n8 VDD.n7 0.00380159
R389 VDD.n25 VDD.n24 0.00380159
R390 VDD.n24 VDD.n23 0.00380159
R391 VDD.n41 VDD.n40 0.00380159
R392 VDD.n40 VDD.n39 0.00380159
R393 VDD.n57 VDD.n56 0.00380159
R394 VDD.n56 VDD.n55 0.00380159
R395 VDD.n74 VDD.n73 0.00380159
R396 VDD.n153 VDD.n152 0.00380159
R397 VDD.n152 VDD.n151 0.00380159
R398 VDD.n183 VDD.n179 0.00380159
R399 VDD.n179 VDD.n178 0.00380159
R400 VDD.n171 VDD.n170 0.00380159
R401 VDD.n170 VDD.n169 0.00380159
R402 VDD.n73 VDD.n72 0.00369982
R403 VDD.n184 VDD.n183 0.00233287
R404 VDD.n172 VDD.n171 0.00233287
R405 VDD.n72 VDD.n71 0.00160176
R406 VDD.n10 VDD.n9 0.000567328
R407 VDD.n26 VDD.n25 0.000567328
R408 VDD.n42 VDD.n41 0.000567328
R409 VDD.n58 VDD.n57 0.000567328
R410 VDD.n75 VDD.n74 0.000567328
R411 VDD.n154 VDD.n153 0.000567328
R412 VDD.n138 VDD.n137 0.000567328
R413 VDD.n122 VDD.n121 0.000567328
R414 VDD.n106 VDD.n105 0.000567328
R415 VDD.n90 VDD.n89 0.000567328
R416 EN.n0 EN.t1 155.304
R417 EN.n0 EN.t0 140.912
R418 EN EN.n0 0.178234
C0 x3.Vin CLK 0.00525f
C1 x4.Vin x2.Vin 1.29e-19
C2 x7.Vin VDD 1.18f
C3 EN a_1696_1902# 0.0121f
C4 x9.Vin CLK 5e-19
C5 x9.Vin x5.Vin 9.41e-20
C6 x11.Vin x2.Vin 0.0031f
C7 x8.Vin x6.Vin 9.41e-20
C8 EN VDD 0.221f
C9 x3.Vin x2.Vin 0.18f
C10 x4.Vin VDD 0.633f
C11 x5.Vin CLK 2.81e-19
C12 x8.Vin x7.Vin 0.18f
C13 x11.Vin VDD 0.628f
C14 x9.Vout VDD 0.633f
C15 x8.Vin VDD 0.636f
C16 x6.Vin x5.Vin 0.184f
C17 x9.Vout x4.Vin 9.79e-20
C18 CLK x2.Vin 0.313f
C19 x3.Vin VDD 0.634f
C20 x5.Vin x2.Vin 5.75e-20
C21 x9.Vin VDD 0.633f
C22 a_1696_1902# CLK 0.0403f
C23 x9.Vout x11.Vin 0.184f
C24 x4.Vin x3.Vin 0.184f
C25 x9.Vin x4.Vin 0.0031f
C26 x6.Vin x2.Vin 1.23e-20
C27 x11.Vin x3.Vin 9.79e-20
C28 x9.Vout x3.Vin 0.0031f
C29 CLK VDD 0.565f
C30 x9.Vout x9.Vin 0.184f
C31 x5.Vin VDD 0.633f
C32 a_1696_1902# x2.Vin 0.1f
C33 x7.Vin x6.Vin 0.177f
C34 x8.Vin x9.Vin 0.184f
C35 EN CLK 0.0385f
C36 x4.Vin CLK 6.89e-19
C37 x5.Vin x4.Vin 0.184f
C38 x6.Vin VDD 0.629f
C39 x11.Vin CLK 0.177f
C40 x9.Vout CLK 0.00103f
C41 x2.Vin VDD 0.853f
C42 x8.Vin CLK 8.14e-20
C43 a_1696_1902# VDD 0.00661f
C44 x8.Vin x5.Vin 0.0031f
C45 EN x2.Vin 0.0787f
C46 EN 0 0.406f
C47 x8.Vin 0 0.583f
C48 x9.Vin 0 0.582f
C49 x9.Vout 0 0.582f
C50 x11.Vin 0 0.597f
C51 a_1696_1902# 0 0.377f $ **FLOATING
C52 x7.Vin 0 0.853f
C53 x6.Vin 0 0.597f
C54 x5.Vin 0 0.582f
C55 x4.Vin 0 0.582f
C56 x3.Vin 0 0.583f
C57 CLK 0 1.15f
C58 x2.Vin 0 0.725f
C59 VDD 0 12.2f
.ends

